[
  {
    "legtypes": [
      {
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            46,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -102,
            63,
            72,
            2,
            81,
            28,
            -57,
            111,
            49,
            105,
            -86,
            92,
            108,
            118,
            -120,
            104,
            58,
            40,
            117,
            -88,
            -31,
            26,
            4,
            65,
            34,
            5,
            -83,
            16,
            3,
            -99,
            -54,
            -91,
            63,
            72,
            81,
            45,
            89,
            32,
            -102,
            -117,
            26,
            104,
            -48,
            31,
            40,
            18,
            42,
            17,
            116,
            -118,
            -122,
            64,
            -109,
            -10,
            -74,
            -38,
            -54,
            -87,
            -75,
            -106,
            -26,
            23,
            -17,
            42,
            -45,
            83,
            59,
            -17,
            -68,
            -13,
            -82,
            -25,
            -17,
            11,
            95,
            -34,
            -32,
            -61,
            -17,
            -17,
            125,
            -18,
            -25,
            79,
            -60,
            71,
            81,
            32,
            16,
            8,
            4,
            2,
            -127,
            64,
            32,
            -114,
            -110,
            -111,
            101,
            -22,
            96,
            111,
            -69,
            -29,
            78,
            70,
            105,
            -91,
            15,
            -2,
            70,
            -91,
            34,
            72,
            113,
            43,
            38,
            53,
            28,
            30,
            91,
            -79,
            78,
            80,
            13,
            -128,
            112,
            16,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            -24,
            82,
            0,
            -50,
            -76,
            -89,
            -128,
            -18,
            -76,
            72,
            -76,
            75,
            26,
            111,
            119,
            3,
            96,
            -83,
            -119,
            19,
            7,
            -32,
            53,
            -85,
            67,
            -121,
            43,
            -26,
            -90,
            -58,
            -81,
            87,
            -10,
            23,
            -75,
            47,
            -126,
            -49,
            63,
            116,
            113,
            -124,
            -44,
            96,
            71,
            102,
            -19,
            -95,
            17,
            -128,
            77,
            -105,
            -107,
            -41,
            -9,
            9,
            67,
            101,
            -65,
            96,
            0,
            83,
            -41,
            89,
            -92,
            6,
            79,
            -25,
            -94,
            -49,
            98,
            1,
            -20,
            -5,
            -57,
            -69,
            27,
            0,
            -74,
            -24,
            57,
            64,
            28,
            0,
            -95,
            115,
            -128,
            20,
            0,
            -43,
            115,
            64,
            80,
            23,
            -112,
            2,
            -96,
            122,
            14,
            8,
            -22,
            2,
            82,
            0,
            -120,
            -2,
            54,
            32,
            9,
            64,
            -51,
            44,
            40,
            104,
            -24,
            -18,
            6,
            -48,
            -22,
            28,
            32,
            23,
            64,
            -117,
            93,
            64,
            52,
            -128,
            -106,
            -70,
            -128,
            -88,
            31,
            67,
            -11,
            6,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            -128,
            52,
            0,
            122,
            -30,
            -69,
            72,
            -65,
            19,
            64,
            -122,
            117,
            63,
            -69,
            118,
            26,
            -64,
            -57,
            77,
            47,
            122,
            58,
            -45,
            -95,
            82,
            98,
            -112,
            93,
            59,
            6,
            -64,
            50,
            99,
            67,
            -13,
            -116,
            -71,
            -95,
            29,
            -74,
            73,
            52,
            16,
            -38,
            -112,
            21,
            64,
            -56,
            55,
            -46,
            52,
            127,
            -43,
            78,
            -93,
            -14,
            101,
            -97,
            124,
            0,
            -16,
            -31,
            -102,
            -123,
            -1,
            120,
            -42,
            50,
            33,
            27,
            0,
            124,
            56,
            -66,
            -4,
            5,
            -21,
            -88,
            124,
            0,
            -8,
            -62,
            -85,
            59,
            65,
            14,
            0,
            -83,
            -26,
            -29,
            78,
            -112,
            28,
            0,
            -29,
            -74,
            -41,
            -124,
            44,
            57,
            109,
            -24,
            42,
            21,
            67,
            -73,
            -103,
            52,
            -54,
            29,
            -89,
            36,
            -123,
            -32,
            58,
            -9,
            20,
            -71,
            -59,
            -57,
            22,
            -121,
            5,
            -27,
            55,
            -126,
            -48,
            22,
            0,
            110,
            0,
            14,
            -82,
            -10,
            -106,
            111,
            -82,
            110,
            -113,
            -108,
            0,
            -60,
            -28,
            11,
            7,
            -64,
            94,
            -108,
            10,
            7,
            -71,
            5,
            -23,
            -125,
            1,
            -34,
            2,
            -80,
            -27,
            2,
            -16,
            120,
            -86,
            19,
            -107,
            -1,
            -5,
            30,
            61,
            -19,
            -3,
            -39,
            -22,
            97,
            -58,
            24,
            81,
            0,
            36,
            -110,
            -46,
            -7,
            -84,
            68,
            125,
            4,
            8,
            -54,
            -57,
            5,
            -28,
            -71,
            67,
            40,
            29,
            -113,
            -80,
            -31,
            -7,
            -109,
            -6,
            33,
            -28,
            97,
            -52,
            101,
            -110,
            -14,
            27,
            62,
            -123,
            102,
            -106,
            37,
            92,
            5,
            -7,
            -108,
            -101,
            49,
            -46,
            -4,
            -31,
            -90,
            119,
            -71,
            -18,
            111,
            40,
            -99,
            -1,
            -3,
            20,
            76,
            -59,
            -65,
            -56,
            -29,
            34,
            73,
            -50,
            -81,
            -56,
            -53,
            -48,
            -3,
            95,
            -45,
            -39,
            -24,
            -59,
            107,
            -89,
            111,
            -13,
            40,
            -99,
            15,
            2,
            -127,
            64,
            32,
            16,
            8,
            -12,
            -81,
            -11,
            9,
            -41,
            90,
            -78,
            9,
            32,
            28,
            68,
            120,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 120.0,
              "Max": 120.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 1000.0,
              "Max": 1000.0
            },
            "id": "#-1:-1",
            "name": "Transportation",
            "lastUpdate": 0,
            "uniqueIdentifier": "adde4589-2e0a-405f-997e-eaf7571b5412",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Truck",
        "lastUpdate": 1448100270026,
        "uniqueIdentifier": "125f1f53-749d-4c83-ad73-467f8e43597c",
        "description": "Truck Transportation"
      },
      {
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            3,
            12,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            -65,
            -117,
            19,
            65,
            20,
            -57,
            -9,
            79,
            -72,
            -54,
            90,
            43,
            -69,
            -13,
            -80,
            -80,
            -112,
            -88,
            -121,
            54,
            106,
            101,
            -93,
            -40,
            8,
            -121,
            88,
            26,
            60,
            -19,
            36,
            -115,
            88,
            8,
            7,
            7,
            -15,
            20,
            20,
            65,
            -16,
            -64,
            31,
            112,
            104,
            97,
            41,
            57,
            97,
            115,
            32,
            22,
            91,
            92,
            -82,
            57,
            11,
            33,
            -39,
            66,
            27,
            109,
            34,
            36,
            7,
            -55,
            -18,
            -31,
            115,
            -65,
            -109,
            -84,
            110,
            -42,
            -51,
            -19,
            36,
            59,
            -69,
            59,
            -77,
            -103,
            7,
            -33,
            38,
            -13,
            118,
            -26,
            -67,
            -49,
            -18,
            -68,
            121,
            -69,
            49,
            12,
            109,
            -38,
            -76,
            105,
            -53,
            -40,
            -18,
            94,
            62,
            79,
            -66,
            52,
            -128,
            89,
            -79,
            -102,
            77,
            11,
            -77,
            13,
            -96,
            -27,
            -42,
            103,
            22,
            -64,
            102,
            -53,
            53,
            -57,
            1,
            -88,
            -75,
            -100,
            70,
            -79,
            -109,
            111,
            -70,
            -9,
            60,
            0,
            52,
            14,
            0,
            -58,
            10,
            -101,
            -68,
            105,
            -45,
            97,
            36,
            24,
            7,
            -128,
            -115,
            -37,
            -5,
            75,
            69,
            75,
            126,
            14,
            -113,
            55,
            47,
            -128,
            -62,
            61,
            9,
            -63,
            -60,
            120,
            1,
            20,
            -94,
            30,
            12,
            -17,
            -68,
            61,
            13,
            0,
            -26,
            -41,
            116,
            94,
            40,
            95,
            -15,
            -61,
            73,
            77,
            2,
            64,
            -23,
            122,
            -16,
            -47,
            -34,
            -65,
            20,
            -107,
            -48,
            -92,
            0,
            6,
            16,
            -2,
            53,
            78,
            42,
            -35,
            -3,
            -74,
            48,
            0,
            -34,
            54,
            -62,
            118,
            82,
            -89,
            -45,
            -13,
            -10,
            -18,
            -72,
            100,
            -90,
            1,
            -96,
            -44,
            -55,
            -128,
            61,
            27,
            -105,
            -56,
            -76,
            0,
            54,
            -101,
            -50,
            -78,
            -12,
            85,
            63,
            54,
            -119,
            36,
            0,
            6,
            106,
            75,
            -35,
            -26,
            102,
            0,
            -128,
            -11,
            8,
            -46,
            -43,
            4,
            -34,
            -32,
            69,
            0,
            -112,
            -86,
            71,
            8,
            -73,
            -71,
            89,
            1,
            -112,
            -90,
            71,
            -120,
            -85,
            -8,
            105,
            2,
            -56,
            -3,
            100,
            64,
            -125,
            50,
            77,
            -48,
            34,
            1,
            -28,
            90,
            15,
            -94,
            -6,
            -4,
            -84,
            1,
            12,
            101,
            74,
            93,
            -11,
            51,
            0,
            -112,
            109,
            61,
            56,
            -88,
            -49,
            -49,
            11,
            0,
            -109,
            -19,
            46,
            74,
            -45,
            -20,
            -28,
            2,
            -64,
            83,
            -86,
            -11,
            -128,
            -89,
            -51,
            -51,
            27,
            64,
            -86,
            61,
            -126,
            -80,
            0,
            83,
            6,
            -112,
            -39,
            -15,
            -120,
            -105,
            19,
            -17,
            36,
            -40,
            -111,
            17,
            64,
            -90,
            -17,
            12,
            -84,
            46,
            12,
            78,
            -123,
            -9,
            18,
            1,
            -96,
            -36,
            -33,
            23,
            88,
            -93,
            20,
            -15,
            -108,
            -120,
            109,
            -124,
            -36,
            58,
            -60,
            -32,
            -29,
            38,
            48,
            57,
            -53,
            56,
            17,
            -92,
            -6,
            -110,
            20,
            124,
            74,
            -8,
            -66,
            10,
            71,
            36,
            -26,
            37,
            37,
            93,
            98,
            73,
            77,
            -1,
            61,
            -82,
            18,
            0,
            42,
            25,
            -90,
            104,
            -19,
            -98,
            59,
            -44,
            -16,
            -107,
            -58,
            -4,
            65,
            37,
            7,
            112,
            -54,
            32,
            69,
            -11,
            -117,
            22,
            -115,
            -71,
            -39,
            5,
            80,
            50,
            -60,
            -68,
            35,
            -48,
            -37,
            53,
            82,
            78,
            -113,
            -17,
            116,
            -60,
            -43,
            0,
            -43,
            -110,
            127,
            -75,
            -14,
            -101,
            110,
            28,
            -97,
            23,
            91,
            8,
            31,
            92,
            -33,
            -91,
            106,
            -103,
            84,
            80,
            122,
            -89,
            -127,
            26,
            123,
            127,
            61,
            -35,
            35,
            -47,
            91,
            64,
            -30,
            -94,
            -73,
            -109,
            106,
            -14,
            15,
            -83,
            -98,
            89,
            -75,
            -100,
            -123,
            56,
            8,
            63,
            -81,
            30,
            -93,
            119,
            111,
            106,
            92,
            65,
            111,
            87,
            -54,
            76,
            60,
            -66,
            -104,
            19,
            115,
            71,
            -114,
            -97,
            52,
            -2,
            -74,
            -55,
            -120,
            17,
            -79,
            -90,
            0,
            -96,
            79,
            -98,
            -38,
            113,
            -37,
            -31,
            -23,
            -42,
            15,
            -8,
            113,
            37,
            53,
            -100,
            -109,
            -37,
            23,
            115,
            71,
            -99,
            -9,
            -95,
            56,
            -37,
            -16,
            77,
            -100,
            -16,
            35,
            -53,
            61,
            -77,
            102,
            -11,
            110,
            -7,
            65,
            -114,
            -54,
            -87,
            126,
            45,
            95,
            -7,
            -32,
            7,
            -15,
            125,
            -23,
            52,
            109,
            -83,
            -82,
            82,
            -108,
            111,
            -93,
            114,
            -109,
            -115,
            -5,
            -66,
            95,
            110,
            95,
            -93,
            -24,
            57,
            -5,
            108,
            44,
            56,
            39,
            -82,
            -115,
            -14,
            -61,
            90,
            108,
            -50,
            97,
            -93,
            -125,
            88,
            17,
            83,
            -108,
            47,
            114,
            -64,
            -8,
            68,
            -55,
            87,
            -83,
            94,
            125,
            92,
            -112,
            -86,
            10,
            57,
            105,
            0,
            26,
            64,
            2,
            0,
            71,
            -98,
            116,
            -24,
            -30,
            70,
            55,
            118,
            33,
            -8,
            -64,
            -105,
            39,
            -88,
            -93,
            -49,
            58,
            76,
            60,
            -66,
            73,
            -41,
            -97,
            10,
            -64,
            -3,
            79,
            125,
            -102,
            127,
            -34,
            97,
            19,
            -6,
            66,
            -64,
            -107,
            122,
            -17,
            -65,
            5,
            -16,
            27,
            -58,
            -126,
            -66,
            -72,
            22,
            115,
            4,
            -3,
            86,
            62,
            -9,
            -87,
            -12,
            -78,
            59,
            -30,
            7,
            -31,
            55,
            -116,
            5,
            125,
            69,
            -82,
            63,
            17,
            -128,
            11,
            27,
            123,
            -33,
            -62,
            11,
            -121,
            -123,
            -59,
            16,
            52,
            20,
            94,
            56,
            44,
            -52,
            -27,
            -5,
            30,
            -28,
            -25,
            -125,
            -128,
            68,
            -81,
            -113,
            -100,
            -72,
            1,
            -100,
            88,
            -17,
            -74,
            -29,
            2,
            85,
            77,
            -56,
            73,
            3,
            -48,
            0,
            52,
            0,
            62,
            59,
            -5,
            122,
            111,
            27,
            23,
            20,
            73,
            -56,
            -55,
            -48,
            -90,
            77,
            -101,
            54,
            109,
            -93,
            -10,
            7,
            -2,
            -101,
            -82,
            76,
            -93,
            53,
            27,
            34,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 120.0,
              "Max": 120.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 1000.0,
              "Max": 1000.0
            },
            "id": "#-1:-1",
            "name": "Transportation",
            "lastUpdate": 0,
            "uniqueIdentifier": "4e856668-3d43-4be0-a791-485592848847",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Barge",
        "lastUpdate": 1448100307814,
        "uniqueIdentifier": "7ce64a22-331d-4a98-8cb1-42febe39fb64",
        "description": "Barge Transportation"
      },
      {
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            3,
            -113,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            93,
            72,
            83,
            97,
            24,
            -57,
            -49,
            -123,
            125,
            -48,
            85,
            87,
            69,
            23,
            97,
            74,
            121,
            25,
            -103,
            20,
            -106,
            19,
            37,
            11,
            -60,
            74,
            103,
            -27,
            -4,
            34,
            -80,
            8,
            2,
            -93,
            24,
            88,
            20,
            89,
            32,
            26,
            73,
            23,
            54,
            3,
            -13,
            99,
            -51,
            102,
            -60,
            10,
            35,
            -102,
            21,
            -107,
            77,
            -99,
            91,
            110,
            -61,
            -87,
            116,
            -68,
            -119,
            46,
            118,
            -31,
            69,
            23,
            125,
            -62,
            81,
            -100,
            -18,
            -104,
            -48,
            -37,
            -98,
            99,
            -109,
            -77,
            -19,
            -52,
            115,
            118,
            60,
            -109,
            109,
            61,
            127,
            -8,
            -63,
            56,
            -25,
            57,
            -49,
            -5,
            60,
            -1,
            -9,
            61,
            -17,
            57,
            71,
            41,
            10,
            -123,
            66,
            -95,
            80,
            40,
            20,
            10,
            -123,
            18,
            -108,
            121,
            -104,
            -34,
            -4,
            -54,
            -22,
            -54,
            19,
            35,
            105,
            13,
            -24,
            -77,
            58,
            -104,
            62,
            -85,
            -109,
            -120,
            50,
            -28,
            52,
            38,
            -87,
            1,
            18,
            -102,
            -1,
            71,
            82,
            27,
            -48,
            -94,
            127,
            68,
            50,
            -10,
            102,
            115,
            8,
            53,
            111,
            -74,
            58,
            38,
            -109,
            -41,
            -128,
            -95,
            -107,
            13,
            48,
            91,
            -99,
            125,
            -80,
            87,
            -4,
            -73,
            43,
            32,
            -87,
            -97,
            2,
            114,
            -18,
            125,
            -46,
            65,
            -39,
            72,
            39,
            69,
            -126,
            104,
            -38,
            52,
            73,
            -54,
            -45,
            73,
            24,
            63,
            115,
            -62,
            25,
            -15,
            -57,
            -38,
            55,
            -112,
            16,
            108,
            104,
            0,
            26,
            -112,
            32,
            123,
            0,
            26,
            -112,
            -116,
            6,
            60,
            125,
            51,
            -64,
            -103,
            0,
            -120,
            26,
            48,
            -80,
            -50,
            68,
            6,
            -41,
            -45,
            -63,
            108,
            -76,
            16,
            107,
            22,
            29,
            70,
            119,
            -54,
            36,
            121,
            -104,
            66,
            7,
            113,
            125,
            -117,
            -123,
            92,
            -35,
            74,
            7,
            113,
            121,
            -101,
            105,
            -51,
            -102,
            110,
            41,
            86,
            25,
            -102,
            -44,
            5,
            -61,
            64,
            -73,
            -18,
            -18,
            -108,
            24,
            -122,
            -94,
            -52,
            -44,
            32,
            3,
            -4,
            -77,
            21,
            54,
            -125,
            48,
            -85,
            66,
            -77,
            29,
            -70,
            82,
            -128,
            -22,
            -44,
            -16,
            -43,
            -94,
            73,
            -29,
            86,
            64,
            -96,
            -82,
            104,
            105,
            59,
            122,
            64,
            43,
            -39,
            -128,
            -38,
            -109,
            106,
            -26,
            72,
            -43,
            57,
            34,
            -107,
            -48,
            -28,
            -79,
            52,
            32,
            -102,
            -70,
            -8,
            -124,
            78,
            -110,
            -94,
            6,
            84,
            106,
            42,
            22,
            -7,
            3,
            -60,
            -54,
            -128,
            -82,
            -62,
            44,
            -107,
            -100,
            -26,
            43,
            -4,
            -11,
            69,
            117,
            11,
            68,
            107,
            0,
            112,
            -19,
            68,
            -95,
            39,
            -106,
            6,
            76,
            -105,
            -19,
            26,
            61,
            91,
            118,
            106,
            94,
            -114,
            1,
            -83,
            -57,
            115,
            -102,
            99,
            110,
            0,
            80,
            82,
            113,
            -6,
            15,
            -36,
            111,
            31,
            -18,
            -19,
            -76,
            -71,
            13,
            -23,
            30,
            62,
            -82,
            -82,
            -116,
            9,
            119,
            -1,
            97,
            79,
            24,
            13,
            -37,
            -61,
            112,
            85,
            101,
            78,
            -72,
            -53,
            -78,
            60,
            -128,
            65,
            83,
            -64,
            -44,
            107,
            -118,
            89,
            -71,
            75,
            -65,
            -13,
            88,
            118,
            121,
            -44,
            -101,
            -96,
            92,
            3,
            -30,
            17,
            89,
            79,
            -127,
            100,
            49,
            -96,
            81,
            125,
            72,
            -2,
            -69,
            -125,
            -81,
            -74,
            84,
            -27,
            -67,
            121,
            -95,
            -97,
            -47,
            -21,
            73,
            34,
            50,
            95,
            87,
            -35,
            -84,
            -56,
            59,
            -63,
            108,
            99,
            -35,
            -89,
            68,
            52,
            64,
            -15,
            -105,
            -93,
            68,
            106,
            126,
            -74,
            65,
            -21,
            81,
            -36,
            0,
            -110,
            67,
            105,
            73,
            -82,
            -1,
            17,
            21,
            -1,
            76,
            -109,
            124,
            42,
            54,
            127,
            -99,
            -126,
            -60,
            -15,
            110,
            64,
            -52,
            -65,
            19,
            -48,
            -128,
            92,
            -86,
            38,
            110,
            13,
            56,
            72,
            -19,
            89,
            -109,
            -81,
            -59,
            120,
            -67,
            -9,
            -41,
            -20,
            115,
            -103,
            -37,
            104,
            -30,
            -51,
            0,
            21,
            -43,
            16,
            -45,
            -90,
            117,
            -29,
            -117,
            -7,
            60,
            3,
            -44,
            43,
            21,
            -13,
            -27,
            76,
            -98,
            -92,
            -94,
            103,
            74,
            118,
            112,
            72,
            -119,
            21,
            -55,
            -87,
            -114,
            84,
            -85,
            98,
            106,
            29,
            91,
            96,
            116,
            -29,
            -84,
            86,
            108,
            21,
            124,
            -84,
            -65,
            72,
            58,
            -20,
            -33,
            37,
            53,
            101,
            50,
            -113,
            113,
            72,
            -119,
            -123,
            -100,
            -112,
            91,
            108,
            -29,
            -125,
            26,
            -95,
            86,
            37,
            27,
            55,
            -6,
            33,
            60,
            -24,
            72,
            -101,
            33,
            52,
            -61,
            -113,
            -75,
            -36,
            127,
            32,
            88,
            -16,
            -24,
            -83,
            27,
            92,
            67,
            -127,
            56,
            -8,
            13,
            -57,
            -124,
            98,
            33,
            7,
            63,
            -89,
            -128,
            97,
            61,
            -68,
            90,
            -23,
            -112,
            90,
            -27,
            -3,
            -61,
            86,
            55,
            -10,
            -69,
            -122,
            107,
            -36,
            -51,
            78,
            -123,
            36,
            12,
            -64,
            -76,
            -37,
            127,
            -67,
            127,
            -85,
            55,
            -39,
            0,
            -45,
            -117,
            -15,
            -49,
            109,
            -50,
            25,
            -97,
            80,
            108,
            -89,
            -19,
            27,
            -13,
            -84,
            119,
            -104,
            14,
            -60,
            26,
            6,
            -89,
            -66,
            70,
            -56,
            73,
            -32,
            92,
            32,
            14,
            -82,
            -127,
            107,
            -123,
            -30,
            96,
            44,
            24,
            19,
            -30,
            58,
            70,
            126,
            52,
            -73,
            -70,
            23,
            -52,
            80,
            -109,
            96,
            -34,
            -91,
            30,
            -116,
            -48,
            83,
            20,
            6,
            -80,
            -74,
            72,
            69,
            38,
            42,
            -48,
            19,
            26,
            -80,
            26,
            3,
            -10,
            25,
            -67,
            -92,
            -34,
            -58,
            -118,
            14,
            4,
            49,
            16,
            43,
            -91,
            -88,
            114,
            -13,
            60,
            -121,
            -108,
            -40,
            -43,
            -114,
            47,
            -37,
            -128,
            75,
            22,
            31,
            -39,
            109,
            -104,
            37,
            105,
            -19,
            75,
            84,
            -66,
            -116,
            92,
            48,
            -100,
            11,
            -60,
            -63,
            53,
            112,
            -83,
            80,
            92,
            -93,
            99,
            -127,
            -88,
            30,
            123,
            -105,
            99,
            11,
            -98,
            -52,
            113,
            -57,
            -124,
            98,
            -107,
            26,
            63,
            42,
            3,
            110,
            -69,
            88,
            -57,
            -107,
            33,
            -106,
            -108,
            62,
            -97,
            91,
            78,
            -56,
            -89,
            -88,
            -41,
            75,
            -50,
            -65,
            99,
            -71,
            -94,
            1,
            -8,
            13,
            -57,
            -124,
            98,
            33,
            7,
            -28,
            -70,
            -29,
            90,
            -102,
            -99,
            -102,
            -41,
            62,
            -63,
            56,
            0,
            -50,
            65,
            12,
            -60,
            42,
            61,
            62,
            -12,
            36,
            -39,
            -128,
            -3,
            61,
            94,
            38,
            82,
            -111,
            -119,
            10,
            -12,
            -124,
            6,
            -96,
            1,
            104,
            0,
            26,
            -128,
            66,
            -95,
            80,
            40,
            20,
            10,
            -123,
            66,
            -95,
            80,
            -96,
            -65,
            63,
            -43,
            -118,
            77,
            -26,
            -69,
            -80,
            -112,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 120.0,
              "Max": 120.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 1000.0,
              "Max": 1000.0
            },
            "id": "#-1:-1",
            "name": "Transportation",
            "lastUpdate": 0,
            "uniqueIdentifier": "f4ca125f-2c9c-4240-b548-88b50a5c7fea",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Cargo Ship",
        "lastUpdate": 1448100337242,
        "uniqueIdentifier": "5de0a31b-2dbd-42ab-af86-6244add4a685",
        "description": "Cargo Ship Transportation"
      },
      {
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            3,
            40,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            49,
            104,
            19,
            81,
            24,
            -57,
            95,
            18,
            115,
            89,
            -69,
            -22,
            98,
            20,
            -36,
            -125,
            56,
            56,
            8,
            102,
            72,
            22,
            29,
            -38,
            49,
            -55,
            -110,
            -93,
            57,
            59,
            -24,
            80,
            5,
            -107,
            6,
            -108,
            28,
            -70,
            40,
            5,
            19,
            -79,
            -112,
            38,
            -90,
            -92,
            4,
            106,
            81,
            20,
            11,
            34,
            72,
            -123,
            -34,
            -91,
            86,
            112,
            -53,
            -71,
            72,
            55,
            11,
            78,
            78,
            73,
            113,
            116,
            120,
            -66,
            119,
            -105,
            11,
            -41,
            -8,
            114,
            -9,
            -102,
            92,
            -102,
            123,
            -71,
            -9,
            -121,
            -1,
            -44,
            -68,
            -21,
            -9,
            -3,
            -18,
            -67,
            -17,
            125,
            -17,
            29,
            0,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            92,
            30,
            20,
            44,
            -125,
            40,
            -84,
            -126,
            -85,
            -80,
            2,
            10,
            112,
            21,
            -44,
            -111,
            21,
            100,
            72,
            116,
            21,
            -60,
            -40,
            76,
            18,
            5,
            -114,
            18,
            -52,
            -38,
            38,
            71,
            105,
            118,
            -110,
            -82,
            -125,
            -103,
            -18,
            91,
            29,
            57,
            105,
            38,
            0,
            -96,
            -32,
            -118,
            -56,
            45,
            55,
            -109,
            101,
            2,
            64,
            119,
            -35,
            -62,
            19,
            113,
            25,
            -88,
            94,
            4,
            48,
            106,
            82,
            7,
            56,
            49,
            -117,
            -27,
            70,
            -2,
            34,
            44,
            -33,
            -65,
            12,
            -17,
            -34,
            -68,
            -114,
            -1,
            30,
            -57,
            -53,
            -55,
            -53,
            85,
            92,
            -19,
            79,
            -22,
            -5,
            -109,
            -45,
            -70,
            -73,
            -27,
            11,
            56,
            1,
            -39,
            -30,
            -72,
            110,
            -121,
            106,
            -98,
            -52,
            72,
            -48,
            52,
            -109,
            85,
            127,
            -44,
            4,
            -58,
            6,
            -64,
            102,
            42,
            -74,
            -3,
            14,
            0,
            79,
            85,
            -111,
            117,
            0,
            -119,
            -108,
            20,
            79,
            102,
            114,
            -117,
            118,
            0,
            58,
            14,
            69,
            -87,
            -51,
            42,
            0,
            35,
            121,
            -121,
            49,
            -92,
            -126,
            53,
            -114,
            125,
            -42,
            -69,
            0,
            42,
            96,
            -114,
            98,
            107,
            82,
            38,
            13,
            -96,
            23,
            -53,
            75,
            -28,
            102,
            -28,
            127,
            87,
            -127,
            70,
            -118,
            -107,
            102,
            6,
            68,
            -57,
            -35,
            109,
            65,
            5,
            68,
            -9,
            -98,
            -99,
            -125,
            -38,
            -117,
            51,
            -16,
            79,
            13,
            5,
            -5,
            6,
            92,
            25,
            26,
            64,
            35,
            -32,
            4,
            0,
            -5,
            -89,
            -71,
            -83,
            38,
            -45,
            -110,
            -22,
            8,
            -99,
            -78,
            57,
            -119,
            15,
            28,
            -65,
            43,
            -52,
            -62,
            -90,
            80,
            -128,
            -86,
            -48,
            34,
            6,
            -121,
            -67,
            25,
            28,
            26,
            -24,
            -111,
            56,
            62,
            11,
            52,
            0,
            122,
            -1,
            35,
            -111,
            -111,
            100,
            119,
            0,
            -12,
            77,
            45,
            -40,
            12,
            103,
            -111,
            -117,
            3,
            19,
            -18,
            55,
            14,
            -36,
            -6,
            -68,
            26,
            -8,
            11,
            95,
            7,
            -85,
            -74,
            113,
            109,
            6,
            -34,
            -23,
            -65,
            -77,
            -114,
            27,
            -12,
            124,
            2,
            0,
            60,
            11,
            -36,
            1,
            -16,
            42,
            -96,
            80,
            39,
            -22,
            -28,
            97,
            -37,
            -29,
            -9,
            33,
            -5,
            -25,
            -110,
            0,
            -96,
            78,
            83,
            47,
            -124,
            104,
            25,
            56,
            -75,
            -82,
            -21,
            71,
            6,
            54,
            2,
            42,
            -36,
            22,
            126,
            -71,
            -106,
            52,
            -55,
            27,
            65,
            -25,
            -92,
            113,
            -63,
            -61,
            75,
            -121,
            -26,
            121,
            100,
            0,
            -86,
            -71,
            12,
            -20,
            1,
            84,
            -64,
            -19,
            -18,
            -128,
            67,
            87,
            -33,
            -74,
            -109,
            119,
            -48,
            -78,
            120,
            27,
            50,
            10,
            -37,
            90,
            55,
            -24,
            -11,
            -128,
            -111,
            -76,
            -45,
            27,
            63,
            14,
            0,
            52,
            11,
            104,
            14,
            48,
            -121,
            39,
            -106,
            -8,
            56,
            76,
            0,
            -80,
            -1,
            -4,
            60,
            20,
            31,
            46,
            -21,
            118,
            6,
            -16,
            49,
            -76,
            -31,
            111,
            0,
            104,
            -81,
            -10,
            53,
            0,
            29,
            -126,
            26,
            57,
            -104,
            74,
            0,
            15,
            -106,
            -27,
            -29,
            117,
            93,
            77,
            65,
            102,
            14,
            -58,
            -88,
            69,
            -48,
            30,
            72,
            -72,
            -60,
            40,
            0,
            -103,
            106,
            27,
            -92,
            -19,
            -25,
            81,
            -53,
            59,
            -121,
            -38,
            93,
            -115,
            25,
            0,
            104,
            123,
            119,
            13,
            -128,
            45,
            -100,
            -35,
            -80,
            -88,
            -49,
            18,
            85,
            -24,
            120,
            9,
            64,
            -17,
            72,
            -20,
            -44,
            9,
            -70,
            10,
            67,
            1,
            51,
            6,
            16,
            84,
            71,
            -102,
            17,
            117,
            -126,
            0,
            58,
            -44,
            -121,
            -95,
            -119,
            -36,
            28,
            127,
            57,
            21,
            -41,
            -115,
            64,
            -3,
            -2,
            116,
            -10,
            -37,
            -113,
            15,
            -105,
            90,
            46,
            1,
            -48,
            -84,
            87,
            -26,
            84,
            -57,
            -31,
            73,
            -21,
            94,
            -79,
            26,
            91,
            42,
            -43,
            -96,
            -23,
            -57,
            43,
            -91,
            22,
            -74,
            49,
            -117,
            40,
            -35,
            0,
            41,
            -46,
            -73,
            2,
            38,
            0,
            96,
            45,
            21,
            -21,
            81,
            43,
            4,
            108,
            55,
            -81,
            -30,
            -104,
            -8,
            118,
            -32,
            54,
            0,
            -86,
            59,
            65,
            111,
            -51,
            -126,
            53,
            17,
            39,
            126,
            -25,
            -23,
            -54,
            -34,
            -20,
            -62,
            -30,
            -66,
            25,
            60,
            42,
            100,
            -123,
            -31,
            -34,
            -2,
            -115,
            24,
            115,
            95,
            -109,
            -82,
            101,
            111,
            -27,
            -83,
            23,
            -88,
            61,
            8,
            105,
            73,
            1,
            -45,
            -82,
            120,
            74,
            -116,
            38,
            50,
            -71,
            54,
            9,
            -128,
            -31,
            121,
            113,
            -86,
            1,
            -104,
            123,
            54,
            -10,
            66,
            -2,
            17,
            -36,
            -38,
            -7,
            -86,
            -37,
            2,
            -95,
            -27,
            111,
            0,
            -23,
            -100,
            54,
            -3,
            75,
            32,
            45,
            117,
            124,
            -69,
            4,
            -116,
            -54,
            61,
            47,
            18,
            -117,
            96,
            70,
            -38,
            2,
            126,
            -111,
            113,
            -128,
            -55,
            105,
            -106,
            -28,
            101,
            -64,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            -59,
            53,
            -94,
            -2,
            1,
            -30,
            75,
            -4,
            -15,
            102,
            86,
            12,
            -80,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 120.0,
              "Max": 120.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 1000.0,
              "Max": 1000.0
            },
            "id": "#-1:-1",
            "name": "Transportation",
            "lastUpdate": 0,
            "uniqueIdentifier": "1d1634c8-2f11-462e-a569-a03b4c379eea",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Plane",
        "lastUpdate": 1448100371322,
        "uniqueIdentifier": "a05af681-5b5e-4de0-8516-fe3b0612b1a7",
        "description": "Plane Transportation"
      },
      {
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            -20,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -102,
            -49,
            107,
            19,
            65,
            20,
            -57,
            -9,
            46,
            -126,
            8,
            10,
            -34,
            -6,
            71,
            72,
            -109,
            102,
            67,
            -110,
            -74,
            -46,
            -60,
            104,
            118,
            87,
            108,
            15,
            10,
            -106,
            122,
            16,
            -107,
            -6,
            -93,
            -121,
            122,
            105,
            -93,
            -26,
            86,
            76,
            53,
            -83,
            -24,
            -55,
            30,
            26,
            60,
            -119,
            85,
            19,
            15,
            -126,
            -126,
            -121,
            120,
            16,
            68,
            -44,
            -69,
            94,
            60,
            -117,
            -121,
            -28,
            63,
            24,
            -9,
            45,
            -99,
            -51,
            -20,
            38,
            -39,
            110,
            -10,
            -57,
            -52,
            36,
            -66,
            7,
            95,
            26,
            102,
            38,
            -17,
            125,
            -33,
            103,
            102,
            118,
            9,
            84,
            81,
            48,
            48,
            48,
            48,
            56,
            71,
            -94,
            -106,
            110,
            39,
            107,
            105,
            -62,
            10,
            -58,
            -2,
            -117,
            -26,
            -109,
            53,
            -75,
            -18,
            110,
            -34,
            -42,
            35,
            117,
            119,
            -68,
            -101,
            -33,
            74,
            -25,
            -40,
            -122,
            119,
            62,
            -86,
            -106,
            28,
            16,
            -52,
            53,
            99,
            124,
            -12,
            -43,
            38,
            109,
            -12,
            -45,
            -113,
            20,
            33,
            127,
            85,
            75,
            -83,
            -17,
            41,
            -26,
            42,
            -88,
            -51,
            -79,
            -33,
            125,
            -38,
            -72,
            91,
            35,
            127,
            10,
            74,
            111,
            -50,
            101,
            65,
            103,
            27,
            -58,
            125,
            -73,
            102,
            -97,
            23,
            118,
            -3,
            2,
            -128,
            -75,
            125,
            114,
            -36,
            -90,
            -7,
            -27,
            105,
            -72,
            97,
            24,
            103,
            26,
            -58,
            111,
            -45,
            28,
            57,
            72,
            -89,
            -9,
            74,
            118,
            -125,
            -17,
            -66,
            -12,
            54,
            15,
            99,
            116,
            -66,
            -8,
            90,
            35,
            126,
            114,
            66,
            109,
            -16,
            32,
            12,
            -128,
            31,
            -109,
            -84,
            -44,
            39,
            89,
            -85,
            -63,
            83,
            79,
            85,
            -14,
            -21,
            103,
            -73,
            121,
            -8,
            12,
            99,
            48,
            7,
            107,
            -122,
            -51,
            -53,
            -67,
            -15,
            66,
            -61,
            -104,
            24,
            -42,
            36,
            -43,
            -64,
            87,
            -32,
            -66,
            -126,
            -26,
            5,
            79,
            60,
            119,
            -66,
            29,
            -44,
            -88,
            23,
            -124,
            48,
            57,
            -31,
            58,
            72,
            123,
            -12,
            -5,
            61,
            15,
            102,
            -22,
            121,
            -110,
            122,
            -100,
            -79,
            4,
            -97,
            97,
            44,
            108,
            -34,
            -111,
            1,
            16,
            -105,
            -124,
            1,
            56,
            -86,
            31,
            35,
            -121,
            102,
            14,
            15,
            45,
            -6,
            -3,
            32,
            -33,
            -123,
            -102,
            82,
            0,
            8,
            -38,
            124,
            88,
            0,
            -3,
            32,
            8,
            1,
            16,
            -44,
            124,
            20,
            0,
            -40,
            28,
            8,
            0,
            1,
            32,
            0,
            4,
            -128,
            0,
            16,
            0,
            2,
            -32,
            15,
            -32,
            -8,
            -62,
            9,
            97,
            0,
            -96,
            -74,
            112,
            0,
            -119,
            -121,
            -86,
            48,
            0,
            80,
            27,
            127,
            12,
            33,
            0,
            4,
            -128,
            0,
            16,
            0,
            2,
            64,
            0,
            8,
            0,
            1,
            -120,
            4,
            48,
            -67,
            -82,
            -109,
            -20,
            -86,
            110,
            -3,
            -115,
            -69,
            73,
            -81,
            90,
            -36,
            1,
            36,
            -14,
            -6,
            64,
            21,
            95,
            68,
            -41,
            52,
            -28,
            -14,
            -86,
            37,
            4,
            -64,
            -20,
            -122,
            -18,
            105,
            42,
            115,
            43,
            -70,
            -45,
            -112,
            -71,
            -23,
            93,
            11,
            -68,
            112,
            5,
            48,
            -67,
            -26,
            52,
            -16,
            -7,
            -21,
            31,
            91,
            -71,
            -7,
            11,
            -10,
            -8,
            -44,
            124,
            120,
            8,
            83,
            -25,
            -69,
            117,
            32,
            55,
            91,
            -117,
            -11,
            0,
            -98,
            -8,
            -3,
            -77,
            67,
            73,
            -77,
            11,
            95,
            89,
            -69,
            -25,
            48,
            -11,
            108,
            -17,
            -67,
            -45,
            -40,
            122,
            56,
            -79,
            -71,
            118,
            94,
            125,
            112,
            -44,
            -126,
            -38,
            116,
            46,
            89,
            -30,
            8,
            96,
            -48,
            -18,
            83,
            93,
            -68,
            122,
            -57,
            -13,
            -56,
            6,
            17,
            -28,
            -20,
            87,
            -117,
            93,
            35,
            4,
            -64,
            -53,
            -73,
            -33,
            122,
            76,
            25,
            -117,
            -53,
            -111,
            3,
            48,
            22,
            111,
            -12,
            -44,
            -127,
            -38,
            66,
            0,
            76,
            -50,
            105,
            3,
            -97,
            1,
            96,
            -108,
            -114,
            -69,
            -41,
            5,
            17,
            -101,
            -61,
            13,
            -63,
            -67,
            -114,
            -13,
            9,
            -48,
            14,
            52,
            62,
            57,
            -89,
            71,
            0,
            -64,
            15,
            72,
            77,
            -36,
            21,
            -16,
            50,
            30,
            -43,
            -15,
            -9,
            -101,
            75,
            24,
            0,
            -70,
            67,
            -42,
            -82,
            71,
            124,
            -9,
            29,
            117,
            92,
            -75,
            -92,
            1,
            32,
            -117,
            16,
            0,
            2,
            -32,
            -10,
            26,
            -44,
            59,
            -78,
            53,
            15,
            -98,
            20,
            -98,
            97,
            -66,
            122,
            -74,
            -27,
            1,
            -96,
            109,
            43,
            34,
            -30,
            100,
            -63,
            -56,
            -79,
            42,
            94,
            94,
            46,
            47,
            -84,
            -108,
            9,
            72,
            -69,
            -74,
            90,
            119,
            -49,
            7,
            21,
            -28,
            -94,
            121,
            -13,
            -105,
            -82,
            -81,
            -72,
            -25,
            21,
            89,
            98,
            -23,
            -18,
            38,
            -95,
            26,
            -91,
            -36,
            -47,
            24,
            -84,
            108,
            29,
            -23,
            -102,
            -84,
            -74,
            -94,
            7,
            80,
            109,
            -39,
            -7,
            -51,
            90,
            -110,
            53,
            -65,
            49,
            -63,
            -20,
            80,
            51,
            -58,
            19,
            -42,
            -36,
            -81,
            -47,
            -122,
            -102,
            -14,
            0,
            40,
            111,
            -42,
            -69,
            -69,
            19,
            -97,
            49,
            7,
            104,
            -77,
            -90,
            124,
            119,
            -65,
            92,
            -19,
            -60,
            15,
            -69,
            -38,
            -111,
            -22,
            89,
            -80,
            84,
            126,
            96,
            48,
            -69,
            82,
            -31,
            112,
            -38,
            42,
            76,
            -67,
            -100,
            -126,
            -127,
            -127,
            -127,
            17,
            34,
            -2,
            1,
            110,
            78,
            -91,
            33,
            7,
            -111,
            -34,
            -72,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 120.0,
              "Max": 120.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 1000.0,
              "Max": 1000.0
            },
            "id": "#-1:-1",
            "name": "Transportation",
            "lastUpdate": 0,
            "uniqueIdentifier": "ddf27b2e-734a-4925-af02-83e1ceaebe85",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Train",
        "lastUpdate": 1448101484262,
        "uniqueIdentifier": "17faea36-e419-4ac9-80ab-fbdbbe77c198",
        "description": "Train Transportation"
      }
    ],
    "categories": [
      {
        "id": null,
        "name": "Costs not accounted",
        "lastUpdate": 1448096669391,
        "uniqueIdentifier": "-1",
        "description": "Default procedure"
      },
      {
        "id": null,
        "name": "CheckUp",
        "lastUpdate": 1448100494972,
        "uniqueIdentifier": "1c112fda-752c-49d8-b50d-6b123555b295",
        "description": "CheckUp of Transport Vehicle"
      },
      {
        "id": null,
        "name": "Unload",
        "lastUpdate": 1448100505208,
        "uniqueIdentifier": "46263709-9590-403d-a6fa-d539dfb72279",
        "description": "Unload"
      },
      {
        "id": null,
        "name": "Load",
        "lastUpdate": 1448100513298,
        "uniqueIdentifier": "8db7d300-65dc-4637-a5a9-db24662c9e65",
        "description": "Load"
      }
    ],
    "events": [
      {
        "dependency": null,
        "probability": {
          "inputValues": [
            {
              "Name": "Mean",
              "Value": {
                "Name": "Mean",
                "Value": 0.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Standard Deviation",
              "Value": {
                "Name": "Standard Deviation",
                "Value": 50.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Lower Bound",
              "Value": {
                "Name": "Lower Bound",
                "Value": 0.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Upper Bound",
              "Value": {
                "Name": "Upper Bound",
                "Value": 1.0E9,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            }
          ],
          "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.NormalDistribution"
        },
        "executionState": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 1000000.0,
              "Max": 1000000.0
            },
            "time": {
              "Min": 26.0,
              "Max": 26.0
            },
            "timeType": "WEEKS",
            "cotwo": {
              "Min": 0.0,
              "Max": 0.0
            },
            "id": "#-1:-1",
            "name": "Embargo Delay",
            "lastUpdate": 0,
            "uniqueIdentifier": "7d1f48c0-9fe4-4cee-b174-ed59ce30f117",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Embargo",
        "lastUpdate": 1448100818373,
        "uniqueIdentifier": "de0c9d05-beac-4890-a10a-42df872e9c27",
        "description": "Embargo"
      },
      {
        "dependency": null,
        "probability": {
          "inputValues": [
            {
              "Name": "Mean",
              "Value": {
                "Name": "Mean",
                "Value": 0.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Standard Deviation",
              "Value": {
                "Name": "Standard Deviation",
                "Value": 20.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Lower Bound",
              "Value": {
                "Name": "Lower Bound",
                "Value": 10.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Upper Bound",
              "Value": {
                "Name": "Upper Bound",
                "Value": 100.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            }
          ],
          "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.NormalDistribution"
        },
        "executionState": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 2.0,
              "Max": 2.0
            },
            "timeType": "WEEKS",
            "cotwo": {
              "Min": 0.0,
              "Max": 0.0
            },
            "id": "#-1:-1",
            "name": "Safety Delay",
            "lastUpdate": 0,
            "uniqueIdentifier": "dbd5c77a-d727-4274-9034-34454ac7d028",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Natural Crisis",
        "lastUpdate": 1448100952648,
        "uniqueIdentifier": "ef78bf1d-d168-43bb-86cd-6ed7582d2834",
        "description": "Earthquake, Tsunami, Hurricane"
      },
      {
        "dependency": null,
        "probability": {
          "inputValues": [
            {
              "Name": "Mean",
              "Value": {
                "Name": "Mean",
                "Value": 0.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Standard Deviation",
              "Value": {
                "Name": "Standard Deviation",
                "Value": 0.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Lower Bound",
              "Value": {
                "Name": "Lower Bound",
                "Value": 50000.0,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            },
            {
              "Name": "Upper Bound",
              "Value": {
                "Name": "Upper Bound",
                "Value": 1.0E9,
                "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.input.DoubleInputValue"
              }
            }
          ],
          "propType": "nl.fontys.sofa.limo.domain.component.event.distribution.NormalDistribution"
        },
        "executionState": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 50000.0,
              "Max": 50000.0
            },
            "time": {
              "Min": 26.0,
              "Max": 26.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 0.0,
              "Max": 0.0
            },
            "id": "#-1:-1",
            "name": "Safety Delay",
            "lastUpdate": 0,
            "uniqueIdentifier": "103fdc1d-46ba-49ee-8d39-7c491a899e40",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "War",
        "lastUpdate": 1448101064318,
        "uniqueIdentifier": "58998e22-077e-4acd-8a12-02e4472e37e5",
        "description": ""
      }
    ],
    "hubtypes": [],
    "hubs": [
      {
        "location": {
          "continent": "Europe",
          "country": {
            "isoNumber3": 250,
            "name": "France",
            "isoAlpha2": "FR",
            "isoAlpha3": "FRA"
          },
          "state": null,
          "town": "Paris",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            90,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -102,
            65,
            78,
            -62,
            64,
            20,
            -122,
            57,
            2,
            55,
            -112,
            35,
            -72,
            81,
            92,
            -104,
            -120,
            27,
            -107,
            13,
            52,
            10,
            -122,
            8,
            36,
            -40,
            106,
            -36,
            0,
            -23,
            -50,
            -96,
            9,
            65,
            99,
            98,
            -94,
            24,
            73,
            -68,
            0,
            55,
            -112,
            27,
            -56,
            9,
            -44,
            -115,
            107,
            -68,
            1,
            -98,
            -128,
            58,
            -81,
            -92,
            -79,
            -116,
            -45,
            98,
            -79,
            13,
            -45,
            121,
            -17,
            37,
            -1,
            -126,
            -66,
            97,
            -24,
            124,
            125,
            51,
            -13,
            -26,
            -47,
            68,
            -126,
            -116,
            -116,
            -116,
            108,
            73,
            86,
            -55,
            -84,
            107,
            32,
            -60,
            0,
            -46,
            61,
            16,
            90,
            0,
            -43,
            76,
            -38,
            2,
            17,
            0,
            2,
            -128,
            -48,
            90,
            7,
            59,
            -38,
            -23,
            -18,
            -26,
            11,
            -24,
            -68,
            -80,
            -101,
            -57,
            53,
            -8,
            -30,
            -98,
            37,
            18,
            1,
            64,
            50,
            -17,
            7,
            -50,
            -36,
            -25,
            -59,
            114,
            -126,
            103,
            52,
            11,
            -97,
            -105,
            8,
            0,
            2,
            0,
            -90,
            15,
            0,
            19,
            -59,
            58,
            -16,
            -48,
            52,
            44,
            -48,
            -19,
            89,
            -59,
            -106,
            -13,
            25,
            -51,
            46,
            -32,
            12,
            -8,
            -6,
            -72,
            104,
            -117,
            0,
            96,
            5,
            -48,
            46,
            -25,
            108,
            17,
            0,
            -84,
            0,
            32,
            -5,
            -69,
            56,
            -52,
            -30,
            6,
            0,
            34,
            0,
            -104,
            0,
            -36,
            -41,
            79,
            50,
            94,
            0,
            -64,
            -121,
            -32,
            -23,
            -21,
            29,
            47,
            0,
            -32,
            83,
            30,
            64,
            -73,
            105,
            -68,
            121,
            1,
            0,
            31,
            -102,
            -7,
            47,
            -114,
            0,
            4,
            -21,
            0,
            1,
            -64,
            12,
            -32,
            -50,
            -84,
            -83,
            -50,
            3,
            0,
            109,
            -108,
            27,
            56,
            -4,
            -3,
            53,
            -81,
            16,
            34,
            40,
            -113,
            105,
            4,
            64,
            -87,
            -71,
            -33,
            -48,
            77,
            119,
            -88,
            -77,
            -49,
            67,
            -105,
            111,
            -56,
            -7,
            -44,
            -85,
            12,
            -15,
            -125,
            100,
            123,
            126,
            -49,
            -107,
            27,
            -12,
            103,
            0,
            52,
            -115,
            -127,
            -46,
            -85,
            63,
            -97,
            -10,
            -70,
            -45,
            99,
            101,
            119,
            -125,
            -103,
            -89,
            -33,
            48,
            62,
            127,
            101,
            -120,
            -20,
            -102,
            -78,
            0,
            -70,
            117,
            67,
            -29,
            -62,
            -65,
            47,
            72,
            -111,
            103,
            -90,
            1,
            124,
            71,
            -119,
            -63,
            63,
            -102,
            -75,
            36,
            31,
            -34,
            -20,
            90,
            74,
            -48,
            46,
            37,
            104,
            -105,
            84,
            111,
            -11,
            -9,
            9,
            111,
            -66,
            29,
            -5,
            110,
            77,
            -71,
            -59,
            47,
            16,
            0,
            21,
            -42,
            2,
            116,
            0,
            74,
            -103,
            -115,
            84,
            117,
            123,
            109,
            11,
            116,
            89,
            -42,
            -6,
            87,
            70,
            -55,
            114,
            -85,
            117,
            -108,
            123,
            114,
            -4,
            -68,
            -64,
            -57,
            -73,
            -121,
            62,
            28,
            63,
            -12,
            45,
            61,
            -128,
            -96,
            41,
            111,
            80,
            17,
            0,
            -39,
            -19,
            -58,
            -40,
            95,
            105,
            21,
            -77,
            19,
            -81,
            -73,
            64,
            22,
            87,
            118,
            2,
            125,
            75,
            15,
            -96,
            93,
            -50,
            127,
            -124,
            63,
            -8,
            -87,
            -38,
            -43,
            -4,
            -85,
            -12,
            0,
            -94,
            26,
            124,
            44,
            -34,
            35,
            -22,
            84,
            11,
            102,
            -44,
            0,
            -32,
            55,
            98,
            -75,
            -25,
            11,
            -78,
            -69,
            119,
            -56,
            -16,
            -32,
            4,
            8,
            -87,
            46,
            -56,
            62,
            13,
            -78,
            107,
            -74,
            -17,
            15,
            125,
            -60,
            22,
            -128,
            -24,
            16,
            52,
            -17,
            80,
            20,
            11,
            0,
            -45,
            3,
            -113,
            62,
            -14,
            123,
            -22,
            11,
            -100,
            33,
            124,
            -94,
            65,
            31,
            73,
            117,
            80,
            98,
            55,
            52,
            -10,
            -70,
            -39,
            -1,
            -36,
            -88,
            -24,
            36,
            -23,
            -126,
            48,
            -114,
            69,
            -24,
            -53,
            -36,
            119,
            56,
            -59,
            14,
            -81,
            57,
            -21,
            42,
            122,
            -122,
            93,
            79,
            12,
            -78,
            -90,
            68,
            106,
            -94,
            90,
            -98,
            95,
            -47,
            99,
            81,
            -29,
            -1,
            80,
            -15,
            -86,
            45,
            74,
            19,
            -6,
            -35,
            -122,
            -15,
            21,
            122,
            -92,
            -79,
            62,
            -91,
            -101,
            10,
            62,
            -85,
            -66,
            25,
            -2,
            111,
            -3,
            -68,
            87,
            -80,
            116,
            0,
            -66,
            -37,
            94,
            -124,
            101,
            44,
            59,
            89,
            -110,
            97,
            91,
            92,
            -26,
            -45,
            -16,
            -39,
            22,
            59,
            9,
            50,
            50,
            50,
            -78,
            -128,
            -10,
            13,
            -120,
            -116,
            43,
            120,
            -15,
            -83,
            113,
            60,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "4e9adb43-71a4-4f4e-af8b-06816479dc45",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "bda2c3ae-fb24-4d44-b2f8-b94ca3af03d1",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Paris",
        "lastUpdate": 1448097197654,
        "uniqueIdentifier": "32cfbd10-626c-4f41-8c60-f2d30da57b58",
        "description": "Paris Logistics Centre"
      },
      {
        "location": {
          "continent": "Europe",
          "country": {
            "isoNumber3": 380,
            "name": "Italy",
            "isoAlpha2": "IT",
            "isoAlpha3": "ITA"
          },
          "state": null,
          "town": "Rome",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            3,
            -51,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            -21,
            75,
            20,
            81,
            24,
            -58,
            -3,
            19,
            -58,
            -11,
            54,
            -21,
            53,
            -95,
            -66,
            68,
            80,
            -87,
            -79,
            88,
            98,
            -117,
            -111,
            38,
            -70,
            90,
            16,
            66,
            10,
            -102,
            -8,
            65,
            36,
            63,
            88,
            40,
            -92,
            -111,
            -122,
            -27,
            37,
            48,
            87,
            -37,
            85,
            49,
            76,
            -117,
            -52,
            34,
            8,
            43,
            100,
            55,
            40,
            88,
            8,
            4,
            -69,
            -48,
            118,
            51,
            34,
            -93,
            -107,
            -120,
            92,
            -115,
            20,
            -22,
            83,
            20,
            -100,
            -10,
            -35,
            -104,
            113,
            -10,
            -20,
            -52,
            56,
            55,
            117,
            118,
            -9,
            60,
            -16,
            -64,
            56,
            -100,
            93,
            124,
            126,
            -25,
            -99,
            115,
            -34,
            51,
            27,
            21,
            69,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            -92,
            76,
            -56,
            117,
            -104,
            66,
            -50,
            -94,
            42,
            -28,
            -80,
            -84,
            68,
            94,
            -8,
            -121,
            -106,
            82,
            -28,
            -76,
            32,
            -42,
            62,
            24,
            -31,
            31,
            -38,
            81,
            60,
            25,
            16,
            58,
            -48,
            -98,
            112,
            15,
            -17,
            22,
            9,
            -49,
            -8,
            120,
            120,
            -123,
            118,
            22,
            -101,
            37,
            -124,
            14,
            112,
            24,
            -123,
            -73,
            -116,
            -55,
            13,
            31,
            22,
            0,
            124,
            -77,
            -18,
            18,
            10,
            -9,
            -5,
            65,
            17,
            -70,
            -45,
            -108,
            -119,
            70,
            -21,
            119,
            -7,
            13,
            -41,
            112,
            47,
            96,
            -100,
            -93,
            -72,
            47,
            108,
            103,
            -100,
            9,
            -114,
            59,
            104,
            -84,
            -93,
            -88,
            33,
            20,
            1,
            32,
            -51,
            0,
            -124,
            -30,
            -114,
            -64,
            13,
            48,
            63,
            118,
            -64,
            111,
            21,
            0,
            2,
            -42,
            -126,
            -71,
            -117,
            113,
            53,
            115,
            -99,
            113,
            93,
            111,
            -37,
            99,
            92,
            -72,
            23,
            7,
            -24,
            -74,
            37,
            59,
            93,
            -11,
            125,
            -112,
            -34,
            -81,
            11,
            0,
            16,
            -100,
            9,
            -74,
            48,
            126,
            80,
            49,
            -128,
            -39,
            14,
            -38,
            -21,
            110,
            53,
            -4,
            122,
            -38,
            28,
            -115,
            -60,
            -20,
            -23,
            -119,
            71,
            94,
            -69,
            -111,
            107,
            -73,
            -41,
            102,
            -100,
            -12,
            -38,
            19,
            74,
            23,
            -122,
            -24,
            45,
            27,
            14,
            -32,
            101,
            127,
            46,
            27,
            12,
            -82,
            -107,
            2,
            -8,
            59,
            85,
            -120,
            -98,
            -73,
            24,
            -48,
            90,
            0,
            -64,
            24,
            0,
            126,
            -37,
            -116,
            43,
            80,
            41,
            43,
            86,
            -118,
            -46,
            21,
            -128,
            -55,
            -106,
            61,
            -126,
            107,
            -122,
            -89,
            111,
            43,
            27,
            -14,
            77,
            123,
            28,
            -21,
            -49,
            -67,
            -23,
            -14,
            1,
            112,
            -68,
            46,
            32,
            -92,
            0,
            -104,
            -71,
            -108,
            -61,
            -69,
            54,
            40,
            -15,
            -46,
            -56,
            78,
            22,
            -64,
            -41,
            126,
            90,
            54,
            -124,
            85,
            -45,
            30,
            77,
            96,
            72,
            1,
            -96,
            -75,
            25,
            0,
            31,
            58,
            98,
            85,
            0,
            -8,
            -1,
            120,
            -88,
            -122,
            -128,
            3,
            -8,
            120,
            37,
            47,
            -72,
            -55,
            -111,
            97,
            -8,
            60,
            -73,
            105,
            114,
            95,
            -50,
            21,
            4,
            96,
            45,
            -93,
            -48,
            41,
            75,
            -70,
            -33,
            -25,
            -54,
            -46,
            -48,
            -93,
            -26,
            36,
            -59,
            48,
            96,
            87,
            81,
            4,
            67,
            -53,
            -103,
            -27,
            86,
            17,
            -41,
            -9,
            -80,
            -11,
            -30,
            -117,
            109,
            27,
            -86,
            51,
            83,
            -24,
            104,
            86,
            52,
            11,
            -128,
            -15,
            -35,
            -122,
            100,
            117,
            85,
            97,
            -89,
            93,
            -78,
            118,
            17,
            -83,
            -62,
            67,
            -43,
            -116,
            -97,
            -52,
            16,
            -36,
            49,
            -96,
            50,
            -104,
            -79,
            -97,
            -122,
            -77,
            -3,
            -31,
            -63,
            45,
            37,
            116,
            0,
            -128,
            -26,
            35,
            105,
            104,
            -34,
            106,
            84,
            -3,
            104,
            104,
            10,
            -32,
            -57,
            -19,
            -126,
            -96,
            64,
            112,
            79,
            -54,
            -20,
            11,
            85,
            -63,
            -43,
            -38,
            116,
            22,
            66,
            83,
            73,
            -102,
            104,
            21,
            -68,
            -18,
            76,
            12,
            -86,
            20,
            -72,
            -89,
            9,
            8,
            41,
            0,
            96,
            -53,
            -61,
            3,
            57,
            -38,
            76,
            -78,
            0,
            -32,
            125,
            -61,
            -30,
            -51,
            -68,
            -43,
            42,
            -80,
            -60,
            -117,
            2,
            -24,
            62,
            -106,
            26,
            4,
            -64,
            90,
            -103,
            42,
            -87,
            26,
            100,
            1,
            120,
            -46,
            -75,
            23,
            -51,
            -12,
            -28,
            40,
            106,
            -123,
            -27,
            2,
            0,
            51,
            0,
            -16,
            -75,
            0,
            7,
            -128,
            -121,
            103,
            -116,
            -121,
            29,
            -83,
            77,
            65,
            19,
            -11,
            41,
            -54,
            0,
            -68,
            27,
            48,
            -77,
            -1,
            40,
            92,
            111,
            4,
            -128,
            10,
            -109,
            118,
            0,
            -90,
            26,
            -109,
            -39,
            -5,
            112,
            45,
            27,
            -128,
            -38,
            86,
            88,
            9,
            -128,
            -23,
            -50,
            12,
            -50,
            98,
            -104,
            -92,
            10,
            0,
            124,
            -122,
            -17,
            -13,
            -70,
            6,
            -64,
            125,
            12,
            -54,
            77,
            84,
            -24,
            3,
            -128,
            -59,
            -46,
            -47,
            106,
            -14,
            27,
            -2,
            102,
            12,
            91,
            32,
            126,
            -62,
            100,
            -36,
            -21,
            107,
            -122,
            -64,
            -89,
            15,
            81,
            -56,
            86,
            17,
            -117,
            -122,
            -85,
            -109,
            -48,
            -83,
            -70,
            4,
            125,
            1,
            88,
            79,
            127,
            27,
            -38,
            46,
            -23,
            -28,
            -8,
            -2,
            -126,
            120,
            -37,
            -84,
            25,
            -128,
            -57,
            -25,
            -77,
            5,
            103,
            107,
            61,
            -4,
            -25,
            126,
            -66,
            36,
            0,
            -81,
            -38,
            12,
            -94,
            0,
            -98,
            -75,
            39,
            -94,
            -63,
            -102,
            20,
            -27,
            0,
            -12,
            -26,
            -97,
            19,
            -39,
            104,
            -7,
            122,
            -90,
            -86,
            -29,
            -13,
            -90,
            1,
            -128,
            -74,
            120,
            118,
            -48,
            -20,
            -85,
            -92,
            -4,
            53,
            -57,
            -62,
            24,
            24,
            43,
            116,
            0,
            123,
            113,
            -42,
            -96,
            31,
            0,
            -16,
            104,
            -120,
            -123,
            -126,
            16,
            124,
            -117,
            37,
            -34,
            54,
            11,
            -75,
            -41,
            96,
            28,
            4,
            -9,
            37,
            10,
            -108,
            57,
            120,
            83,
            0,
            112,
            27,
            37,
            -104,
            49,
            -66,
            49,
            -16,
            -30,
            -124,
            47,
            20,
            -2,
            59,
            2,
            -2,
            59,
            3,
            -41,
            -16,
            29,
            -36,
            -17,
            92,
            -66,
            -106,
            -27,
            15,
            63,
            82,
            73,
            -15,
            54,
            58,
            27,
            2,
            -32,
            70,
            -61,
            110,
            -34,
            80,
            66,
            -128,
            -8,
            12,
            91,
            35,
            51,
            22,
            -82,
            -59,
            -58,
            -30,
            -99,
            40,
            -45,
            49,
            114,
            -49,
            12,
            -16,
            -2,
            64,
            83,
            0,
            -52,
            -84,
            -64,
            -87,
            13,
            47,
            67,
            -83,
            27,
            -95,
            -75,
            -58,
            -31,
            -37,
            48,
            -45,
            44,
            -99,
            -56,
            -117,
            22,
            -20,
            3,
            -32,
            8,
            13,
            80,
            -70,
            -53,
            83,
            3,
            -114,
            -45,
            -70,
            -20,
            4,
            -107,
            2,
            -64,
            -49,
            12,
            33,
            -37,
            10,
            -53,
            5,
            80,
            -67,
            -113,
            -30,
            61,
            58,
            71,
            12,
            -128,
            -58,
            -126,
            -104,
            -43,
            -105,
            39,
            -123,
            49,
            -111,
            7,
            -64,
            121,
            102,
            7,
            -17,
            99,
            16,
            49,
            0,
            -72,
            111,
            -113,
            52,
            7,
            64,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            68,
            20,
            9,
            -6,
            7,
            -84,
            22,
            112,
            24,
            61,
            -101,
            -52,
            -61,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "1dcaae7d-b0a9-4a0c-980d-9b6c38717b4b",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "9464ff11-44f1-4c51-88fc-4f7c4c4e74b4",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Rome",
        "lastUpdate": 1448097133334,
        "uniqueIdentifier": "732f7bc0-7ee3-4d93-af23-4e257679e035",
        "description": "Rome Logistics Centre"
      },
      {
        "location": {
          "continent": "Europe",
          "country": {
            "isoNumber3": 826,
            "name": "United Kingdom",
            "isoAlpha2": "GB",
            "isoAlpha3": "GBR"
          },
          "state": null,
          "town": "London",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            -117,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -102,
            -49,
            43,
            4,
            97,
            24,
            -57,
            -3,
            9,
            -82,
            -110,
            85,
            44,
            37,
            68,
            14,
            -82,
            28,
            112,
            96,
            -107,
            -93,
            -44,
            30,
            -44,
            30,
            20,
            23,
            46,
            118,
            29,
            52,
            -105,
            89,
            9,
            -75,
            69,
            -111,
            3,
            -79,
            73,
            14,
            123,
            34,
            -78,
            14,
            -42,
            117,
            71,
            -10,
            -64,
            -51,
            -123,
            -125,
            66,
            98,
            -83,
            -108,
            -94,
            125,
            -19,
            51,
            118,
            -58,
            -76,
            59,
            51,
            118,
            -52,
            46,
            -13,
            62,
            -17,
            -5,
            -42,
            -73,
            -90,
            103,
            -26,
            125,
            -89,
            -17,
            -89,
            -9,
            -57,
            51,
            -17,
            59,
            101,
            101,
            -68,
            -4,
            95,
            -15,
            -49,
            72,
            -99,
            32,
            102,
            1,
            4,
            -126,
            82,
            -52,
            31,
            -108,
            -114,
            89,
            6,
            64,
            64,
            -52,
            25,
            23,
            -124,
            68,
            121,
            64,
            -108,
            -98,
            20,
            0,
            112,
            13,
            49,
            118,
            -58,
            -66,
            24,
            15,
            -87,
            -26,
            -77,
            -126,
            24,
            115,
            93,
            63,
            87,
            -52,
            -52,
            -4,
            70,
            0,
            -104,
            88,
            17,
            -116,
            -52,
            51,
            -45,
            11,
            -104,
            5,
            -112,
            55,
            -13,
            27,
            9,
            -21,
            -118,
            -96,
            55,
            -13,
            27,
            -50,
            5,
            24,
            87,
            -124,
            66,
            -51,
            -93,
            28,
            10,
            -28,
            -64,
            35,
            -112,
            -125,
            126,
            98,
            77,
            30,
            -127,
            3,
            -64,
            8,
            64,
            24,
            -86,
            -105,
            -75,
            50,
            -42,
            -92,
            -102,
            93,
            30,
            109,
            86,
            -29,
            -52,
            0,
            -48,
            -102,
            -43,
            -117,
            113,
            0,
            28,
            0,
            18,
            0,
            126,
            81,
            18,
            -84,
            46,
            -127,
            -33,
            -7,
            -128,
            68,
            55,
            -124,
            41,
            49,
            -34,
            -6,
            91,
            -13,
            -118,
            -96,
            13,
            -118,
            83,
            -33,
            120,
            -62,
            46,
            0,
            104,
            -125,
            -54,
            -44,
            -40,
            -74,
            113,
            -102,
            51,
            -61,
            64,
            -16,
            116,
            -96,
            -40,
            0,
            -96,
            77,
            58,
            -52,
            23,
            -93,
            -37,
            -101,
            12,
            7,
            -57,
            3,
            88,
            -101,
            11,
            29,
            -105,
            82,
            -114,
            7,
            112,
            -69,
            84,
            65,
            20,
            93,
            -50,
            127,
            73,
            27,
            3,
            93,
            -52,
            86,
            22,
            20,
            -45,
            -85,
            79,
            13,
            0,
            48,
            52,
            -29,
            117,
            -53,
            -46,
            -102,
            88,
            -12,
            -43,
            -54,
            9,
            -49,
            -55,
            116,
            -107,
            26,
            -117,
            78,
            -71,
            -28,
            -40,
            -22,
            72,
            13,
            -7,
            -87,
            62,
            53,
            0,
            -10,
            38,
            -85,
            -43,
            -20,
            14,
            -82,
            -107,
            -72,
            54,
            -21,
            51,
            -117,
            25,
            -43,
            -25,
            0,
            56,
            0,
            39,
            126,
            -20,
            -20,
            123,
            18,
            -42,
            55,
            60,
            108,
            42,
            -13,
            78,
            7,
            125,
            -19,
            -3,
            -79,
            -7,
            -84,
            28,
            15,
            32,
            -71,
            -47,
            -104,
            -73,
            -76,
            89,
            85,
            42,
            -36,
            66,
            39,
            -128,
            -41,
            -19,
            118,
            -37,
            -26,
            21,
            65,
            91,
            -44,
            1,
            120,
            -39,
            106,
            43,
            26,
            0,
            104,
            11,
            13,
            -128,
            -69,
            -43,
            58,
            66,
            -34,
            -82,
            117,
            5,
            -9,
            -48,
            3,
            72,
            63,
            -97,
            27,
            2,
            -128,
            123,
            104,
            1,
            60,
            108,
            119,
            -28,
            25,
            -34,
            -36,
            9,
            -53,
            -54,
            -115,
            -61,
            -77,
            -24,
            0,
            -68,
            -33,
            28,
            -27,
            25,
            -19,
            30,
            -14,
            -55,
            -54,
            -115,
            -65,
            -33,
            68,
            -15,
            1,
            -48,
            -21,
            -14,
            70,
            0,
            64,
            76,
            0,
            -24,
            -54,
            -104,
            7,
            41,
            67,
            65,
            59,
            28,
            80,
            1,
            120,
            62,
            -12,
            -103,
            -10,
            0,
            -83,
            -108,
            123,
            79,
            -69,
            -125,
            120,
            0,
            60,
            70,
            -6,
            44,
            3,
            -128,
            58,
            -24,
            -121,
            -128,
            -103,
            -48,
            -51,
            1,
            -23,
            -44,
            69,
            -63,
            -26,
            -31,
            89,
            116,
            0,
            82,
            -79,
            -15,
            -126,
            1,
            -64,
            -77,
            40,
            51,
            65,
            -77,
            52,
            -40,
            44,
            29,
            70,
            -107,
            10,
            -61,
            -20,
            110,
            100,
            94,
            59,
            -13,
            -93,
            5,
            -64,
            -4,
            -41,
            32,
            51,
            0,
            62,
            118,
            123,
            -56,
            -3,
            -118,
            -53,
            -74,
            121,
            104,
            3,
            -38,
            -94,
            114,
            75,
            -116,
            -99,
            61,
            -63,
            125,
            -49,
            -43,
            63,
            -20,
            10,
            95,
            57,
            107,
            107,
            60,
            -38,
            -37,
            10,
            -1,
            -11,
            36,
            -41,
            27,
            98,
            -91,
            -108,
            -4,
            -65,
            81,
            -26,
            93,
            84,
            28,
            -114,
            -106,
            66,
            -44,
            -100,
            12,
            -99,
            -119,
            -107,
            -22,
            -55,
            14,
            92,
            43,
            -15,
            -123,
            97,
            -73,
            28,
            -117,
            76,
            124,
            -97,
            -10,
            -64,
            53,
            -60,
            -32,
            -34,
            79,
            -11,
            -47,
            28,
            -115,
            105,
            -51,
            6,
            -67,
            110,
            126,
            54,
            -56,
            1,
            112,
            0,
            72,
            0,
            -16,
            -62,
            11,
            93,
            -27,
            19,
            -69,
            118,
            -4,
            -83,
            77,
            -25,
            86,
            -78,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "69edd686-d912-46f7-8602-fdf78fd2c4fb",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "6e8685f1-1210-4da8-a905-33103dae2ad6",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "London",
        "lastUpdate": 1448097330369,
        "uniqueIdentifier": "52c883ff-9327-4d85-ab1a-c06753778044",
        "description": "London Logistics Centre"
      },
      {
        "location": {
          "continent": "Asia",
          "country": {
            "isoNumber3": 356,
            "name": "India",
            "isoAlpha2": "IN",
            "isoAlpha3": "IND"
          },
          "state": null,
          "town": "Dehli",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            -84,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -104,
            -51,
            74,
            -61,
            64,
            16,
            -57,
            125,
            4,
            31,
            -63,
            71,
            -24,
            27,
            -24,
            -35,
            -117,
            -24,
            73,
            16,
            44,
            8,
            -118,
            8,
            126,
            -32,
            65,
            4,
            -123,
            98,
            65,
            68,
            80,
            20,
            60,
            9,
            18,
            15,
            -94,
            -94,
            -120,
            86,
            60,
            120,
            81,
            11,
            -74,
            -43,
            -74,
            72,
            20,
            -12,
            -96,
            -88,
            -24,
            69,
            18,
            61,
            -12,
            17,
            98,
            -89,
            -72,
            -110,
            -90,
            -101,
            102,
            -109,
            76,
            -46,
            124,
            -52,
            -64,
            -128,
            -44,
            -51,
            -50,
            127,
            126,
            -101,
            -39,
            -39,
            77,
            91,
            27,
            25,
            25,
            25,
            25,
            25,
            25,
            25,
            89,
            11,
            76,
            -38,
            127,
            -47,
            -64,
            9,
            64,
            92,
            109,
            -9,
            -24,
            109,
            22,
            60,
            -74,
            0,
            114,
            37,
            -75,
            2,
            30,
            -53,
            -60,
            -13,
            37,
            85,
            -45,
            123,
            44,
            64,
            -28,
            75,
            -33,
            9,
            99,
            -30,
            -115,
            -2,
            -99,
            -120,
            100,
            -14,
            -123,
            -94,
            -38,
            -61,
            91,
            121,
            -34,
            -101,
            0,
            99,
            -93,
            -74,
            -14,
            73,
            -21,
            -107,
            111,
            120,
            19,
            -110,
            49,
            78,
            62,
            34,
            16,
            -60,
            106,
            62,
            -94,
            123,
            -126,
            44,
            87,
            -38,
            69,
            106,
            94,
            100,
            79,
            -128,
            -71,
            66,
            -72,
            -6,
            110,
            87,
            -66,
            -34,
            67,
            -107,
            -4,
            -115,
            92,
            -23,
            -64,
            6,
            0,
            115,
            6,
            -78,
            -75,
            -15,
            90,
            86,
            -82,
            -84,
            76,
            98,
            3,
            -128,
            57,
            69,
            -29,
            -5,
            82,
            -33,
            85,
            81,
            -110,
            78,
            -96,
            -92,
            -81,
            -45,
            124,
            81,
            61,
            -63,
            6,
            0,
            115,
            -42,
            -59,
            47,
            -86,
            -57,
            102,
            -15,
            -3,
            -88,
            111,
            -103,
            35,
            82,
            -42,
            1,
            72,
            121,
            0,
            32,
            37,
            26,
            -33,
            -29,
            -28,
            -107,
            -84,
            -7,
            -114,
            -83,
            92,
            -71,
            -17,
            -3,
            -51,
            -49,
            4,
            34,
            -15,
            91,
            -70,
            -69,
            -21,
            74,
            4,
            21,
            0,
            123,
            -59,
            91,
            -38,
            45,
            -102,
            -47,
            111,
            124,
            11,
            -16,
            -37,
            -96,
            -99,
            -8,
            94,
            109,
            124,
            -62,
            -85,
            -107,
            47,
            42,
            31,
            120,
            -11,
            -81,
            124,
            -40,
            -115,
            -113,
            -33,
            -37,
            -53,
            63,
            93,
            -62,
            61,
            -69,
            58,
            -10,
            -17,
            -34,
            -65,
            -115,
            112,
            18,
            -36,
            118,
            26,
            31,
            -65,
            4,
            -124,
            -38,
            -101,
            -78,
            -58,
            -5,
            -18,
            -25,
            -44,
            -35,
            -58,
            -9,
            -67,
            12,
            -52,
            62,
            124,
            98,
            0,
            112,
            18,
            -33,
            -77,
            47,
            -71,
            34,
            -126,
            -79,
            1,
            56,
            -119,
            79,
            0,
            -126,
            126,
            -53,
            11,
            -35,
            -83,
            -111,
            0,
            -60,
            5,
            -128,
            -76,
            -9,
            -100,
            -30,
            -43,
            24,
            -106,
            -48,
            -125,
            -45,
            119,
            109,
            96,
            44,
            91,
            115,
            -8,
            27,
            107,
            94,
            -18,
            -34,
            80,
            -51,
            -59,
            83,
            0,
            59,
            -121,
            -81,
            -38,
            -6,
            -26,
            -109,
            -80,
            -56,
            -12,
            -22,
            -3,
            127,
            -14,
            -52,
            -31,
            55,
            -47,
            -25,
            -41,
            54,
            31,
            107,
            49,
            125,
            3,
            -112,
            94,
            41,
            115,
            1,
            100,
            -50,
            63,
            -75,
            -95,
            -87,
            -21,
            -70,
            68,
            -84,
            -60,
            27,
            -57,
            -21,
            29,
            -2,
            103,
            -11,
            -68,
            113,
            60,
            104,
            -32,
            1,
            -48,
            107,
            118,
            5,
            96,
            110,
            -15,
            70,
            75,
            116,
            74,
            92,
            0,
            -68,
            100,
            -74,
            118,
            -97,
            77,
            -59,
            -61,
            -86,
            -103,
            37,
            47,
            82,
            14,
            48,
            -73,
            21,
            52,
            -90,
            19,
            52,
            -125,
            118,
            -41,
            0,
            96,
            34,
            -16,
            -15,
            -39,
            108,
            3,
            0,
            59,
            73,
            -116,
            -50,
            20,
            44,
            -109,
            103,
            14,
            99,
            -101,
            -19,
            25,
            70,
            55,
            2,
            0,
            -83,
            76,
            55,
            26,
            -128,
            -2,
            -31,
            51,
            87,
            0,
            68,
            -109,
            55,
            43,
            37,
            59,
            0,
            122,
            7,
            51,
            -8,
            0,
            -70,
            -5,
            -113,
            28,
            3,
            -128,
            58,
            -75,
            11,
            -64,
            88,
            -37,
            118,
            0,
            -128,
            -42,
            64,
            1,
            -32,
            -43,
            -82,
            -107,
            27,
            -9,
            -110,
            80,
            3,
            -128,
            -74,
            101,
            23,
            0,
            60,
            19,
            8,
            0,
            24,
            7,
            33,
            12,
            0,
            -127,
            62,
            8,
            17,
            -128,
            -72,
            3,
            -104,
            95,
            -70,
            -45,
            102,
            -46,
            101,
            -33,
            0,
            76,
            -52,
            -35,
            -42,
            98,
            -6,
            6,
            -128,
            -99,
            1,
            -116,
            0,
            -106,
            55,
            30,
            44,
            -5,
            55,
            38,
            -128,
            -53,
            -36,
            -105,
            -27,
            56,
            -90,
            -77,
            47,
            -103,
            -63,
            1,
            48,
            50,
            125,
            97,
            122,
            20,
            -26,
            9,
            -25,
            93,
            106,
            -80,
            0,
            44,
            -84,
            -54,
            66,
            93,
            -128,
            117,
            47,
            -48,
            -114,
            -42,
            6,
            -39,
            100,
            97,
            104,
            -125,
            108,
            -47,
            -24,
            28,
            64,
            0,
            8,
            0,
            1,
            112,
            12,
            -128,
            -116,
            -116,
            -116,
            -116,
            -116,
            -116,
            44,
            -14,
            -10,
            11,
            -24,
            70,
            24,
            -93,
            -72,
            66,
            55,
            -113,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "f547e81c-a776-4458-827b-0b482b9b7633",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "92eb1cba-2837-4455-a8ea-61c0bf38773d",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Dehli",
        "lastUpdate": 1448099049520,
        "uniqueIdentifier": "bb89d804-62db-472b-903b-257d8c3c44c6",
        "description": "Dehli Logistics Centre"
      },
      {
        "location": {
          "continent": "NorthAmerica",
          "country": {
            "isoNumber3": 840,
            "name": "United States",
            "isoAlpha2": "US",
            "isoAlpha3": "USA"
          },
          "state": null,
          "town": "Washington DC",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            1,
            -69,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            -65,
            78,
            -61,
            48,
            16,
            -58,
            -5,
            8,
            60,
            2,
            -113,
            -64,
            27,
            -64,
            0,
            123,
            87,
            42,
            -122,
            74,
            116,
            99,
            -23,
            35,
            -28,
            1,
            -112,
            -102,
            25,
            -119,
            102,
            108,
            -38,
            -111,
            25,
            -87,
            8,
            53,
            -96,
            6,
            -119,
            48,
            -80,
            36,
            -107,
            96,
            67,
            4,
            6,
            51,
            -77,
            24,
            95,
            -107,
            -128,
            84,
            -30,
            34,
            74,
            112,
            -3,
            -25,
            59,
            -23,
            -109,
            -94,
            75,
            28,
            -5,
            126,
            113,
            -20,
            -69,
            -92,
            -47,
            -128,
            -63,
            96,
            -80,
            53,
            -39,
            94,
            -85,
            -61,
            73,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            -32,
            -110,
            -19,
            -18,
            119,
            -70,
            101,
            -16,
            -91,
            -56,
            -25,
            18,
            -128,
            -73,
            111,
            0,
            90,
            -121,
            -52,
            25,
            0,
            81,
            -100,
            -13,
            42,
            1,
            0,
            0,
            0,
            0,
            0,
            88,
            111,
            -63,
            32,
            107,
            7,
            97,
            -58,
            43,
            37,
            -50,
            -39,
            15,
            64,
            22,
            124,
            33,
            -85,
            -125,
            -65,
            -66,
            121,
            -35,
            25,
            -98,
            61,
            -68,
            -53,
            -126,
            -89,
            115,
            116,
            -115,
            85,
            65,
            39,
            9,
            -37,
            -104,
            -60,
            -49,
            99,
            -39,
            123,
            47,
            19,
            -75,
            -95,
            -74,
            -58,
            3,
            -104,
            -60,
            57,
            -5,
            109,
            -16,
            95,
            16,
            114,
            115,
            -77,
            -61,
            40,
            126,
            105,
            -81,
            26,
            -8,
            -94,
            -82,
            -90,
            121,
            -45,
            -87,
            39,
            111,
            -4,
            76,
            -120,
            -90,
            -71,
            87,
            87,
            -16,
            -97,
            18,
            -9,
            52,
            99,
            -91,
            79,
            -40,
            102,
            -19,
            -63,
            23,
            -94,
            123,
            59,
            53,
            -11,
            -115,
            124,
            21,
            -2,
            43,
            120,
            99,
            -46,
            101,
            103,
            1,
            -120,
            76,
            -82,
            -9,
            83,
            -102,
            91,
            -93,
            122,
            -102,
            21,
            56,
            -87,
            -89,
            48,
            -8,
            -94,
            112,
            74,
            -11,
            -39,
            21,
            -6,
            97,
            122,
            -89,
            26,
            0,
            -11,
            -87,
            -47,
            -12,
            -97,
            117,
            -107,
            -49,
            0,
            -47,
            -89,
            -42,
            -117,
            -96,
            127,
            114,
            -49,
            15,
            -114,
            46,
            -26,
            -94,
            -29,
            -46,
            95,
            -6,
            72,
            -53,
            124,
            -78,
            -10,
            -58,
            -20,
            2,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            96,
            55,
            -128,
            -2,
            104,
            -74,
            -67,
            -88,
            -13,
            -53,
            39,
            78,
            58,
            29,
            100,
            -36,
            59,
            -66,
            -99,
            -117,
            -114,
            75,
            127,
            -23,
            35,
            45,
            -13,
            -55,
            -38,
            87,
            -11,
            -87,
            62,
            -11,
            29,
            101,
            91,
            65,
            -104,
            62,
            -86,
            79,
            127,
            101,
            18,
            99,
            17,
            99,
            82,
            89,
            -6,
            114,
            29,
            -91,
            18,
            -128,
            -81,
            33,
            0,
            -33,
            -2,
            111,
            0,
            -70,
            125,
            27,
            88,
            101,
            21,
            -1,
            -21,
            46,
            80,
            117,
            -19,
            -38,
            -73,
            60,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            112,
            7,
            64,
            48,
            76,
            -101,
            34,
            3,
            99,
            26,
            -91,
            -63,
            -116,
            -58,
            -92,
            -78,
            22,
            96,
            26,
            -42,
            2,
            76,
            37,
            0,
            -57,
            -85,
            65,
            -99,
            10,
            33,
            29,
            127,
            -106,
            -62,
            96,
            48,
            99,
            -20,
            3,
            63,
            -20,
            -2,
            67,
            54,
            105,
            97,
            -7,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "4b7bf3ab-d724-43a9-b9b2-3618f10b25d7",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "9e59b26b-28e9-449d-ac60-4764f3357c31",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Washington",
        "lastUpdate": 1448099066121,
        "uniqueIdentifier": "fe0b91ba-73e9-4b52-b817-34e9f3fbe072",
        "description": "Washington Logistics Centre"
      },
      {
        "location": {
          "continent": "Europe",
          "country": {
            "isoNumber3": 724,
            "name": "Spain",
            "isoAlpha2": "ES",
            "isoAlpha3": "ESP"
          },
          "state": null,
          "town": "Madrid",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            4,
            -16,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            -49,
            79,
            19,
            65,
            20,
            -57,
            -3,
            19,
            -4,
            19,
            -8,
            19,
            122,
            -127,
            94,
            48,
            46,
            -119,
            18,
            126,
            -87,
            32,
            24,
            68,
            64,
            26,
            64,
            84,
            44,
            -92,
            -32,
            15,
            48,
            64,
            93,
            36,
            -31,
            -105,
            16,
            -118,
            -119,
            -63,
            68,
            12,
            96,
            107,
            -112,
            122,
            -112,
            -77,
            96,
            -38,
            3,
            23,
            -115,
            9,
            28,
            -71,
            -63,
            -63,
            59,
            77,
            76,
            -72,
            -82,
            -13,
            -74,
            -99,
            118,
            -103,
            -50,
            -18,
            -68,
            -74,
            -77,
            -37,
            -42,
            -20,
            36,
            47,
            -30,
            -18,
            -20,
            123,
            -33,
            -7,
            -52,
            -101,
            -97,
            -67,
            116,
            -55,
            45,
            110,
            113,
            -117,
            91,
            36,
            22,
            127,
            -109,
            -94,
            14,
            53,
            -43,
            104,
            105,
            107,
            80,
            124,
            -7,
            -6,
            -126,
            111,
            -115,
            -66,
            -64,
            119,
            -55,
            3,
            -72,
            -48,
            120,
            -35,
            -108,
            -77,
            64,
            -99,
            82,
            -111,
            -85,
            31,
            -8,
            6,
            -66,
            101,
            -3,
            -107,
            33,
            -128,
            -4,
            122,
            46,
            43,
            -109,
            -54,
            25,
            64,
            62,
            -61,
            -128,
            77,
            -1,
            -14,
            1,
            64,
            -124,
            -5,
            27,
            107,
            18,
            84,
            -16,
            96,
            -125,
            -30,
            -55,
            -41,
            23,
            124,
            -101,
            -50,
            34,
            -16,
            89,
            -64,
            124,
            -30,
            104,
            -127,
            -15,
            59,
            59,
            -40,
            -93,
            77,
            118,
            -75,
            -50,
            23,
            -22,
            11,
            124,
            -128,
            -81,
            124,
            -26,
            -111,
            -94,
            -106,
            -83,
            -7,
            87,
            -38,
            -42,
            92,
            112,
            -77,
            96,
            63,
            -60,
            7,
            -8,
            42,
            -69,
            -27,
            48,
            5,
            32,
            46,
            1,
            64,
            -68,
            -20,
            0,
            108,
            44,
            -88,
            -51,
            58,
            0,
            9,
            -62,
            -87,
            31,
            -16,
            89,
            18,
            -115,
            -37,
            -100,
            127,
            117,
            6,
            -126,
            -56,
            -65,
            49,
            81,
            -81,
            -55,
            4,
            -80,
            53,
            31,
            -36,
            -75,
            -48,
            116,
            -104,
            -46,
            116,
            102,
            107,
            -29,
            63,
            45,
            -88,
            -127,
            -116,
            32,
            -46,
            43,
            115,
            106,
            -123,
            9,
            -128,
            83,
            -39,
            0,
            72,
            -29,
            78,
            -72,
            -39,
            70,
            52,
            24,
            53,
            -127,
            70,
            123,
            -46,
            122,
            78,
            85,
            -116,
            -127,
            -52,
            -120,
            -77,
            -11,
            -28,
            101,
            -128,
            14,
            92,
            -55,
            -18,
            -3,
            96,
            -126,
            -43,
            -59,
            -85,
            103,
            19,
            -128,
            96,
            2,
            -111,
            37,
            -118,
            -84,
            -104,
            -97,
            -26,
            84,
            95,
            -47,
            0,
            96,
            -121,
            -128,
            113,
            -4,
            -89,
            86,
            2,
            53,
            -1,
            -34,
            15,
            -122,
            24,
            95,
            -15,
            -94,
            13,
            -127,
            44,
            -30,
            38,
            75,
            92,
            86,
            -113,
            20,
            -80,
            20,
            -78,
            48,
            -51,
            -26,
            1,
            90,
            -113,
            -105,
            -111,
            -46,
            -53,
            -34,
            78,
            88,
            -35,
            -113,
            70,
            -76,
            -40,
            -10,
            118,
            -123,
            104,
            -52,
            22,
            58,
            15,
            96,
            125,
            -127,
            22,
            -48,
            -76,
            -9,
            53,
            18,
            -80,
            31,
            64,
            52,
            -110,
            -128,
            96,
            -5,
            -47,
            112,
            8,
            43,
            -102,
            55,
            118,
            -123,
            -61,
            -115,
            124,
            -125,
            5,
            0,
            90,
            82,
            -102,
            -50,
            108,
            7,
            -112,
            12,
            68,
            104,
            71,
            -61,
            -36,
            -44,
            126,
            122,
            -89,
            -2,
            47,
            107,
            -109,
            -99,
            -73,
            -65,
            -28,
            124,
            6,
            32,
            -33,
            -16,
            124,
            113,
            53,
            -19,
            -124,
            -113,
            -88,
            46,
            -57,
            0,
            -104,
            5,
            -29,
            29,
            97,
            71,
            90,
            -82,
            -97,
            -25,
            26,
            103,
            -92,
            -91,
            -10,
            28,
            123,
            28,
            22,
            105,
            114,
            12,
            -64,
            120,
            103,
            83,
            59,
            -9,
            62,
            32,
            -113,
            115,
            -68,
            -103,
            -97,
            -119,
            -114,
            27,
            -43,
            69,
            3,
            -16,
            61,
            -6,
            -39,
            99,
            21,
            108,
            121,
            -72,
            87,
            93,
            30,
            -18,
            -45,
            120,
            -58,
            -42,
            -19,
            82,
            -68,
            -95,
            110,
            -59,
            -85,
            37,
            -83,
            114,
            37,
            -37,
            23,
            -33,
            15,
            -60,
            -80,
            2,
            0,
            26,
            109,
            3,
            -16,
            35,
            -6,
            -39,
            103,
            12,
            22,
            -5,
            -74,
            113,
            -39,
            -8,
            126,
            105,
            -72,
            47,
            -124,
            1,
            -48,
            -91,
            84,
            -87,
            -103,
            -58,
            39,
            13,
            -98,
            97,
            0,
            64,
            -116,
            11,
            43,
            0,
            -47,
            96,
            -44,
            4,
            26,
            109,
            92,
            1,
            -62,
            113,
            99,
            48,
            88,
            18,
            -103,
            12,
            56,
            -63,
            0,
            96,
            27,
            79,
            13,
            9,
            -32,
            -112,
            -73,
            44,
            -117,
            38,
            103,
            -23,
            -29,
            63,
            25,
            44,
            -78,
            -117,
            75,
            91,
            121,
            0,
            88,
            95,
            -96,
            -127,
            -43,
            -27,
            72,
            -6,
            -13,
            -126,
            89,
            -119,
            94,
            9,
            -8,
            -46,
            -61,
            -59,
            -89,
            120,
            46,
            -109,
            57,
            -32,
            52,
            -109,
            -2,
            -34,
            83,
            120,
            70,
            -33,
            67,
            93,
            44,
            0,
            -98,
            38,
            91,
            -122,
            1,
            -101,
            -2,
            -23,
            44,
            48,
            -20,
            -66,
            -84,
            68,
            47,
            -7,
            -5,
            -78,
            46,
            52,
            120,
            61,
            -81,
            -49,
            37,
            -92,
            46,
            6,
            0,
            -60,
            -26,
            106,
            -78,
            99,
            24,
            100,
            118,
            -128,
            -84,
            101,
            118,
            -124,
            86,
            -94,
            121,
            -77,
            -73,
            25,
            0,
            -85,
            -43,
            -60,
            8,
            96,
            127,
            39,
            -78,
            105,
            -94,
            73,
            -2,
            -114,
            16,
            35,
            -56,
            18,
            -64,
            80,
            111,
            28,
            13,
            -128,
            -44,
            45,
            52,
            94,
            89,
            3,
            -128,
            -103,
            -66,
            -28,
            0,
            -16,
            14,
            38,
            -58,
            3,
            -54,
            27,
            127,
            -65,
            98,
            61,
            4,
            46,
            -118,
            -70,
            -89,
            84,
            -122,
            -70,
            -110,
            19,
            -96,
            6,
            127,
            99,
            97,
            -125,
            65,
            44,
            -116,
            38,
            71,
            1,
            -120,
            38,
            46,
            -80,
            -59,
            -128,
            -49,
            -109,
            90,
            1,
            98,
            -39,
            27,
            33,
            111,
            12,
            -34,
            97,
            64,
            58,
            14,
            -128,
            119,
            29,
            -58,
            6,
            19,
            77,
            92,
            96,
            -3,
            117,
            87,
            14,
            -52,
            -10,
            0,
            -44,
            6,
            -22,
            -81,
            -2,
            18,
            -7,
            -95,
            19,
            -86,
            -107,
            38,
            -87,
            -41,
            98,
            112,
            -83,
            37,
            10,
            38,
            -102,
            -72,
            -64,
            -4,
            55,
            -81,
            -59,
            83,
            -37,
            -34,
            -29,
            110,
            -91,
            -54,
            -48,
            -16,
            -86,
            -44,
            51,
            -81,
            94,
            71,
            8,
            -128,
            -60,
            18,
            117,
            74,
            33,
            87,
            113,
            -62,
            -85,
            41,
            -34,
            -123,
            7,
            6,
            -64,
            -53,
            -50,
            -26,
            -97,
            -92,
            -111,
            1,
            -46,
            -32,
            56,
            -89,
            -9,
            119,
            -31,
            -35,
            -44,
            -3,
            -42,
            35,
            12,
            0,
            -77,
            11,
            19,
            25,
            87,
            113,
            57,
            -115,
            127,
            -6,
            27,
            -96,
            56,
            109,
            51,
            -5,
            120,
            -85,
            -83,
            -80,
            104,
            5,
            -96,
            6,
            63,
            -108,
            -120,
            116,
            -55,
            26,
            -1,
            21,
            -94,
            64,
            -101,
            -77,
            83,
            7,
            24,
            -47,
            116,
            37,
            -80,
            2,
            -128,
            -11,
            3,
            49,
            69,
            -70,
            -52,
            126,
            -72,
            41,
            -24,
            42,
            -36,
            -52,
            -100,
            6,
            -128,
            -47,
            -108,
            -49,
            93,
            100,
            -50,
            19,
            32,
            -75,
            -43,
            103,
            -125,
            -114,
            1,
            -128,
            88,
            24,
            77,
            82,
            38,
            66,
            -47,
            4,
            72,
            -19,
            -19,
            11,
            63,
            10,
            0,
            -39,
            -12,
            120,
            -52,
            0,
            -64,
            59,
            -116,
            -113,
            119,
            99,
            67,
            88,
            0,
            113,
            -57,
            0,
            -84,
            77,
            4,
            80,
            0,
            -70,
            -107,
            74,
            -97,
            25,
            0,
            -78,
            20,
            54,
            99,
            124,
            64,
            44,
            -25,
            0,
            96,
            2,
            17,
            -5,
            -96,
            62,
            71,
            2,
            -32,
            46,
            -127,
            -23,
            -91,
            16,
            -29,
            99,
            125,
            122,
            76,
            -61,
            -22,
            114,
            12,
            -64,
            -6,
            -52,
            75,
            36,
            0,
            -21,
            -99,
            32,
            -58,
            -57,
            71,
            18,
            -85,
            -28,
            0,
            96,
            87,
            2,
            25,
            0,
            114,
            -47,
            -28,
            2,
            112,
            1,
            20,
            25,
            -64,
            72,
            91,
            -125,
            -42,
            87,
            91,
            -83,
            45,
            62,
            -23,
            65,
            3,
            -128,
            -70,
            -16,
            -51,
            104,
            91,
            125,
            -7,
            3,
            -96,
            13,
            27,
            -17,
            -72,
            -123,
            6,
            0,
            117,
            -83,
            50,
            -94,
            100,
            1,
            80,
            -47,
            -77,
            -113,
            -70,
            -77,
            0,
            60,
            110,
            -84,
            65,
            3,
            -128,
            -70,
            44,
            -128,
            -103,
            7,
            -9,
            -46,
            -49,
            74,
            6,
            0,
            -37,
            35,
            84,
            -96,
            -38,
            -37,
            46,
            29,
            0,
            -8,
            100,
            1,
            96,
            50,
            66,
            26,
            0,
            -40,
            126,
            -66,
            -97,
            26,
            45,
            121,
            0,
            -17,
            39,
            71,
            47,
            108,
            -107,
            -91,
            0,
            0,
            -89,
            -68,
            96,
            -91,
            8,
            -128,
            62,
            3,
            -51,
            -46,
            0,
            24,
            -9,
            -7,
            -27,
            2,
            -128,
            -98,
            23,
            92,
            0,
            46,
            0,
            9,
            -57,
            -31,
            -75,
            -119,
            -111,
            -29,
            -43,
            -47,
            -121,
            9,
            48,
            -3,
            120,
            -100,
            50,
            -6,
            108,
            -3,
            -11,
            -72,
            110,
            3,
            117,
            87,
            117,
            -101,
            -18,
            -67,
            -5,
            91,
            -65,
            36,
            37,
            70,
            -97,
            13,
            -33,
            -86,
            -3,
            3,
            -1,
            79,
            -98,
            6,
            -51,
            13,
            -22,
            64,
            93,
            -6,
            29,
            -11,
            3,
            62,
            -23,
            51,
            26,
            -49,
            74,
            19,
            104,
            -106,
            122,
            49,
            -22,
            22,
            -73,
            -72,
            -59,
            45,
            -1,
            99,
            -7,
            7,
            123,
            28,
            10,
            -106,
            76,
            -117,
            92,
            86,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "db153459-dc92-4d9a-a4f7-ed4a7c93cb7b",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "72caf17e-1528-4340-96c6-6c7f262bd82a",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Madrid",
        "lastUpdate": 1448099131876,
        "uniqueIdentifier": "350a84e3-b75f-403e-a60d-973a22f16d21",
        "description": "Madrid Logistics Centre"
      },
      {
        "location": {
          "continent": "NorthAmerica",
          "country": {
            "isoNumber3": 124,
            "name": "Canada",
            "isoAlpha2": "CA",
            "isoAlpha3": "CAN"
          },
          "state": null,
          "town": "Toronto",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            3,
            -86,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            90,
            -35,
            106,
            19,
            65,
            20,
            62,
            -113,
            -48,
            71,
            -24,
            35,
            -12,
            13,
            -52,
            35,
            108,
            65,
            47,
            -12,
            66,
            -126,
            -105,
            34,
            73,
            68,
            65,
            20,
            -91,
            65,
            81,
            -63,
            34,
            6,
            81,
            -101,
            -10,
            38,
            121,
            3,
            -13,
            6,
            -55,
            27,
            -104,
            55,
            -120,
            55,
            109,
            -75,
            8,
            73,
            106,
            -75,
            -74,
            -43,
            -82,
            115,
            118,
            -77,
            -35,
            100,
            50,
            -65,
            -69,
            -99,
            -39,
            -97,
            -50,
            -127,
            67,
            -62,
            102,
            33,
            -7,
            -66,
            57,
            -25,
            59,
            -33,
            -52,
            6,
            -64,
            -123,
            11,
            23,
            46,
            92,
            20,
            47,
            -4,
            45,
            -88,
            -106,
            9,
            -52,
            -86,
            -42,
            -3,
            109,
            -16,
            49,
            -53,
            67,
            64,
            27,
            -66,
            -8,
            29,
            88,
            81,
            -66,
            -73,
            -124,
            4,
            72,
            1,
            -7,
            59,
            -80,
            70,
            -18,
            25,
            71,
            -9,
            -106,
            -122,
            0,
            127,
            27,
            -68,
            11,
            80,
            -28,
            -67,
            -116,
            -92,
            -14,
            17,
            64,
            -83,
            42,
            -35,
            10,
            -28,
            90,
            -121,
            5,
            -66,
            20,
            4,
            16,
            -15,
            -85,
            48,
            -128,
            93,
            -24,
            1,
            -66,
            -14,
            -64,
            -105,
            -125,
            -128,
            54,
            -116,
            68,
            0,
            101,
            89,
            26,
            -15,
            115,
            4,
            92,
            69,
            2,
            -120,
            -30,
            55,
            -46,
            18,
            -96,
            107,
            -96,
            -14,
            103,
            126,
            20,
            -127,
            -98,
            127,
            -48,
            34,
            102,
            -94,
            106,
            -86,
            -116,
            -6,
            112,
            -47,
            61,
            -8,
            -103,
            42,
            -96,
            -109,
            87,
            57,
            108,
            -117,
            89,
            -7,
            85,
            -91,
            -13,
            -99,
            -77,
            18,
            -28,
            -77,
            -98,
            42,
            -96,
            -33,
            -49,
            -76,
            90,
            98,
            96,
            87,
            -68,
            56,
            36,
            -52,
            -51,
            -9,
            -111,
            9,
            -15,
            -53,
            92,
            20,
            69,
            95,
            76,
            -101,
            -101,
            52,
            4,
            40,
            -81,
            -66,
            -83,
            -107,
            -113,
            -74,
            -82,
            -116,
            31,
            80,
            -99,
            3,
            -41,
            23,
            41,
            -11,
            -126,
            -9,
            -105,
            -28,
            -113,
            59,
            -118,
            4,
            -104,
            22,
            61,
            -115,
            -15,
            -43,
            103,
            92,
            91,
            -48,
            -126,
            37,
            -17,
            -49,
            -55,
            -15,
            93,
            -16,
            -113,
            30,
            43,
            -83,
            126,
            -45,
            -10,
            -8,
            106,
            37,
            -104,
            -41,
            85,
            -35,
            -14,
            -33,
            91,
            7,
            -1,
            -17,
            -69,
            28,
            -107,
            126,
            106,
            -1,
            -66,
            13,
            27,
            -94,
            -99,
            29,
            61,
            -9,
            85,
            -6,
            -65,
            -112,
            -10,
            85,
            37,
            15,
            31,
            40,
            -104,
            31,
            -45,
            -91,
            31,
            -120,
            -35,
            14,
            92,
            91,
            -56,
            54,
            -44,
            77,
            -125,
            -57,
            -66,
            -57,
            -14,
            -49,
            92,
            -12,
            102,
            123,
            -15,
            -119,
            -115,
            21,
            -97,
            -49,
            -3,
            27,
            97,
            -26,
            -90,
            -12,
            109,
            -126,
            -57,
            -78,
            -105,
            -119,
            95,
            -74,
            103,
            118,
            -78,
            -47,
            117,
            47,
            -3,
            -22,
            31,
            63,
            23,
            -10,
            125,
            37,
            43,
            -31,
            -21,
            -87,
            -10,
            -17,
            -7,
            -89,
            -28,
            4,
            72,
            122,
            127,
            88,
            -120,
            -61,
            11,
            -84,
            -126,
            -61,
            -121,
            -20,
            -21,
            103,
            111,
            -59,
            -82,
            79,
            -42,
            -5,
            -63,
            24,
            69,
            113,
            14,
            71,
            42,
            109,
            -70,
            122,
            -90,
            -89,
            66,
            87,
            -107,
            0,
            86,
            43,
            -32,
            53,
            94,
            121,
            -29,
            -106,
            23,
            87,
            31,
            -57,
            95,
            -30,
            22,
            18,
            28,
            -87,
            -101,
            62,
            -59,
            93,
            -56,
            127,
            -17,
            9,
            -40,
            90,
            8,
            -8,
            -24,
            9,
            105,
            -119,
            -113,
            -32,
            79,
            -22,
            98,
            2,
            16,
            -68,
            116,
            -12,
            -119,
            61,
            65,
            55,
            87,
            -83,
            -16,
            -25,
            101,
            92,
            9,
            -40,
            14,
            -47,
            -5,
            -109,
            -41,
            -53,
            -9,
            -94,
            -30,
            -89,
            38,
            -64,
            -58,
            -22,
            -21,
            84,
            1,
            -26,
            -12,
            126,
            12,
            28,
            -13,
            -41,
            83,
            -66,
            -23,
            -63,
            -34,
            -105,
            -6,
            126,
            113,
            126,
            -74,
            -3,
            64,
            -29,
            43,
            -21,
            -121,
            32,
            -120,
            -88,
            -36,
            89,
            73,
            -117,
            99,
            -76,
            -14,
            60,
            -37,
            -117,
            -19,
            35,
            19,
            79,
            78,
            -114,
            2,
            -95,
            36,
            -18,
            -43,
            106,
            21,
            -80,
            64,
            -45,
            -124,
            28,
            -65,
            -120,
            15,
            59,
            68,
            -91,
            -113,
            -32,
            -125,
            -10,
            -87,
            -91,
            54,
            88,
            35,
            124,
            -80,
            106,
            -25,
            96,
            68,
            97,
            58,
            96,
            98,
            -55,
            71,
            -32,
            121,
            -62,
            40,
            -46,
            13,
            -99,
            19,
            98,
            115,
            109,
            16,
            62,
            -82,
            86,
            -2,
            49,
            -89,
            -101,
            -15,
            116,
            -120,
            -64,
            127,
            -65,
            25,
            106,
            -59,
            -23,
            -101,
            112,
            122,
            -80,
            8,
            -96,
            -81,
            107,
            29,
            -113,
            -101,
            88,
            121,
            -99,
            83,
            29,
            -90,
            -35,
            -67,
            30,
            19,
            -64,
            -45,
            10,
            97,
            -42,
            -108,
            72,
            25,
            -102,
            28,
            -125,
            -11,
            -76,
            -101,
            29,
            -52,
            111,
            -73,
            -12,
            -128,
            79,
            27,
            68,
            55,
            54,
            -108,
            -66,
            103,
            104,
            100,
            -69,
            28,
            108,
            -113,
            -73,
            96,
            -112,
            20,
            -4,
            -76,
            30,
            -125,
            -105,
            57,
            -66,
            -97,
            -113,
            -8,
            -114,
            50,
            115,
            67,
            -108,
            -12,
            -103,
            94,
            4,
            94,
            -59,
            -16,
            -96,
            103,
            72,
            66,
            64,
            54,
            -101,
            -92,
            -80,
            50,
            -70,
            60,
            111,
            112,
            -74,
            -87,
            -90,
            -6,
            -84,
            -7,
            95,
            8,
            2,
            4,
            62,
            97,
            -120,
            -32,
            -25,
            87,
            -2,
            -32,
            -74,
            58,
            24,
            36,
            42,
            -63,
            -7,
            -62,
            40,
            55,
            36,
            28,
            120,
            -80,
            70,
            64,
            79,
            34,
            -16,
            73,
            -20,
            46,
            -114,
            -57,
            4,
            27,
            -93,
            74,
            94,
            -64,
            47,
            -10,
            125,
            104,
            -100,
            122,
            -42,
            -114,
            -40,
            108,
            62,
            45,
            -102,
            -113,
            125,
            15,
            -86,
            52,
            -8,
            61,
            15,
            90,
            -78,
            125,
            68,
            -54,
            63,
            74,
            12,
            102,
            -39,
            12,
            -38,
            47,
            -85,
            42,
            -40,
            -11,
            -96,
            67,
            -125,
            23,
            -40,
            -24,
            -98,
            -62,
            54,
            -73,
            81,
            -104,
            127,
            124,
            -116,
            61,
            88,
            -95,
            -63,
            -17,
            -82,
            -117,
            29,
            -103,
            -92,
            26,
            90,
            -123,
            1,
            -65,
            84,
            -14,
            104,
            115,
            61,
            -11,
            30,
            100,
            86,
            -125,
            -19,
            -121,
            -98,
            9,
            75,
            126,
            -52,
            -24,
            -9,
            -60,
            110,
            44,
            -24,
            -31,
            34,
            16,
            16,
            -88,
            -68,
            7,
            125,
            -42,
            -54,
            95,
            -38,
            17,
            124,
            94,
            9,
            96,
            -82,
            122,
            -104,
            -105,
            -70,
            -9,
            54,
            -74,
            -107,
            77,
            9,
            -66,
            -55,
            2,
            -113,
            98,
            -89,
            -45,
            -13,
            -123,
            12,
            50,
            -33,
            43,
            -84,
            85,
            39,
            -83,
            -32,
            -63,
            85,
            8,
            66,
            -64,
            106,
            26,
            -91,
            47,
            77,
            -96,
            -54,
            35,
            25,
            -32,
            -62,
            -123,
            11,
            23,
            46,
            -118,
            31,
            -1,
            1,
            -93,
            -99,
            -119,
            -94,
            61,
            30,
            50,
            103,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "86f70acb-d59a-480e-9469-c9ab72f3f28d",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "f9a362ae-da11-4d17-b2d8-4ea393b09351",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Toronto",
        "lastUpdate": 1448099164238,
        "uniqueIdentifier": "3769b7b4-9bdb-4b98-9608-80f8d5a3221c",
        "description": "Toronto Logistics Centre"
      },
      {
        "location": {
          "continent": "Europe",
          "country": {
            "isoNumber3": 276,
            "name": "Germany",
            "isoAlpha2": "DE",
            "isoAlpha3": "DEU"
          },
          "state": null,
          "town": "Berlin",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            1,
            -12,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -104,
            -65,
            74,
            -61,
            80,
            20,
            -58,
            125,
            -124,
            62,
            -126,
            -113,
            -48,
            -51,
            -47,
            -45,
            77,
            -46,
            43,
            116,
            115,
            114,
            114,
            -46,
            -90,
            82,
            80,
            -60,
            41,
            13,
            93,
            90,
            5,
            -87,
            56,
            -120,
            -109,
            -115,
            -40,
            14,
            86,
            -60,
            93,
            42,
            117,
            119,
            -55,
            -28,
            -30,
            -96,
            111,
            -96,
            111,
            16,
            -17,
            -119,
            36,
            -83,
            37,
            -122,
            -124,
            36,
            109,
            -2,
            124,
            31,
            28,
            -72,
            -71,
            -51,
            -67,
            57,
            -25,
            -41,
            123,
            114,
            111,
            -50,
            -54,
            10,
            4,
            65,
            16,
            4,
            45,
            69,
            -115,
            42,
            53,
            -9,
            20,
            42,
            23,
            50,
            120,
            117,
            -109,
            106,
            -86,
            66,
            -113,
            -11,
            42,
            13,
            -102,
            27,
            -76,
            90,
            72,
            8,
            117,
            -123,
            -124,
            42,
            -120,
            10,
            -101,
            2,
            -86,
            -78,
            -2,
            42,
            1,
            88,
            -71,
            14,
            -110,
            -105,
            -73,
            -52,
            -11,
            15,
            -9,
            -70,
            70,
            37,
            59,
            -8,
            106,
            -27,
            -109,
            -125,
            -73,
            77,
            -90,
            -125,
            -45,
            -17,
            -62,
            17,
            52,
            -55,
            77,
            -82,
            55,
            68,
            -59,
            114,
            -14,
            -100,
            -105,
            -68,
            -99,
            -1,
            -126,
            116,
            7,
            -128,
            -4,
            -3,
            -123,
            -81,
            -25,
            -57,
            -28,
            -26,
            5,
            -87,
            -118,
            -118,
            -55,
            1,
            53,
            4,
            125,
            113,
            80,
            118,
            91,
            -82,
            -118,
            -33,
            -66,
            105,
            -37,
            -34,
            25,
            -28,
            61,
            -36,
            -106,
            64,
            -50,
            115,
            18,
            60,
            -111,
            27,
            104,
            72,
            -53,
            -59,
            -18,
            16,
            5,
            64,
            46,
            86,
            -64,
            77,
            -73,
            101,
            69,
            -79,
            116,
            4,
            -47,
            -47,
            -12,
            48,
            78,
            95,
            28,
            -20,
            90,
            103,
            -5,
            59,
            -74,
            69,
            5,
            -32,
            -52,
            -61,
            115,
            -122,
            26,
            43,
            125,
            -114,
            13,
            64,
            -65,
            -89,
            -105,
            -78,
            6,
            -128,
            125,
            -114,
            117,
            21,
            -12,
            79,
            -12,
            -102,
            -47,
            -43,
            -66,
            -45,
            14,
            -128,
            125,
            100,
            95,
            19,
            75,
            7,
            -98,
            60,
            -83,
            0,
            18,
            13,
            124,
            86,
            -114,
            83,
            105,
            -77,
            -123,
            -67,
            20,
            11,
            5,
            -32,
            -7,
            126,
            -40,
            -102,
            -73,
            -21,
            -10,
            -15,
            36,
            -115,
            -26,
            -27,
            107,
            100,
            0,
            -29,
            -47,
            -64,
            -54,
            -78,
            69,
            6,
            -16,
            52,
            26,
            -106,
            -57,
            119,
            -73,
            102,
            -26,
            -126,
            -105,
            62,
            -77,
            -17,
            -79,
            -91,
            66,
            -31,
            -2,
            -7,
            -1,
            -12,
            112,
            -43,
            51,
            29,
            -69,
            108,
            29,
            -67,
            -77,
            121,
            -11,
            25,
            -89,
            -19,
            55,
            -89,
            -113,
            -37,
            126,
            -9,
            -58,
            57,
            126,
            -95,
            59,
            -64,
            54,
            -83,
            -39,
            -26,
            -43,
            119,
            -72,
            37,
            -36,
            62,
            110,
            -5,
            -35,
            27,
            -25,
            120,
            0,
            40,
            -22,
            25,
            0,
            0,
            0,
            96,
            65,
            0,
            -126,
            22,
            48,
            -126,
            -44,
            16,
            2,
            23,
            77,
            102,
            -66,
            -19,
            -105,
            94,
            64,
            -119,
            15,
            -128,
            102,
            78,
            -25,
            -44,
            -52,
            -20,
            0,
            -24,
            104,
            -122,
            -113,
            -93,
            -58,
            -33,
            34,
            -118,
            119,
            96,
            -13,
            -33,
            -20,
            -2,
            -75,
            6,
            -51,
            -100,
            45,
            110,
            4,
            125,
            126,
            -94,
            10,
            115,
            -6,
            10,
            115,
            74,
            -117,
            50,
            103,
            -94,
            -89,
            63,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            40,
            54,
            0,
            8,
            -126,
            32,
            8,
            -126,
            114,
            -95,
            31,
            65,
            -74,
            -17,
            -101,
            -111,
            29,
            49,
            -12,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "b5740306-b264-4243-a5ab-63a27e411c4e",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "14d3e175-ec3f-4514-94ed-25ac73df1d9e",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Berlin",
        "lastUpdate": 1448099188496,
        "uniqueIdentifier": "8e45cc00-0823-4ec0-a0c3-0dd9cd835c9f",
        "description": "Berlin Logistics Centre"
      },
      {
        "location": {
          "continent": "Asia",
          "country": {
            "isoNumber3": 156,
            "name": "China",
            "isoAlpha2": "CN",
            "isoAlpha3": "CHN"
          },
          "state": null,
          "town": "Peking",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            1,
            -35,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            65,
            78,
            -62,
            64,
            20,
            -122,
            103,
            111,
            72,
            88,
            -80,
            35,
            105,
            112,
            -43,
            89,
            122,
            3,
            79,
            64,
            -30,
            13,
            -12,
            6,
            122,
            3,
            -36,
            -69,
            97,
            7,
            106,
            12,
            -36,
            -96,
            120,
            -126,
            118,
            -125,
            46,
            -23,
            -46,
            -72,
            -87,
            71,
            -32,
            6,
            117,
            94,
            83,
            48,
            41,
            109,
            90,
            -37,
            -95,
            125,
            -45,
            -7,
            95,
            -14,
            39,
            4,
            94,
            -104,
            -9,
            127,
            -76,
            -61,
            123,
            83,
            33,
            16,
            8,
            4,
            2,
            -127,
            -24,
            36,
            62,
            -91,
            -100,
            -111,
            -84,
            52,
            -65,
            117,
            -35,
            -51,
            -121,
            -108,
            113,
            34,
            -41,
            -11,
            -84,
            50,
            127,
            52,
            -98,
            17,
            0,
            88,
            4,
            96,
            -99,
            3,
            96,
            109,
            13,
            -128,
            -35,
            100,
            50,
            84,
            123,
            64,
            120,
            48,
            79,
            -81,
            -23,
            61,
            -85,
            -10,
            -127,
            120,
            41,
            124,
            -91,
            56,
            -107,
            111,
            -101,
            -7,
            56,
            79,
            118,
            -104,
            95,
            -120,
            -69,
            34,
            0,
            -12,
            89,
            -65,
            -51,
            63,
            -117,
            89,
            -95,
            -7,
            -125,
            84,
            -114,
            13,
            -9,
            124,
            -103,
            -4,
            62,
            25,
            -113,
            -2,
            97,
            60,
            -85,
            -56,
            100,
            -29,
            -9,
            13,
            -51,
            31,
            33,
            -88,
            -37,
            -30,
            -106,
            -73,
            -39,
            23,
            113,
            69,
            69,
            -86,
            98,
            119,
            26,
            12,
            -105,
            105,
            -105,
            -84,
            -91,
            -42,
            -28,
            -16,
            43,
            -17,
            91,
            48,
            92,
            -90,
            125,
            -73,
            -65,
            -4,
            82,
            -124,
            29,
            -102,
            15,
            89,
            92,
            9,
            9,
            -116,
            -107,
            24,
            -86,
            75,
            -13,
            -26,
            123,
            58,
            14,
            -50,
            41,
            90,
            -125,
            -42,
            50,
            110,
            -46,
            -45,
            37,
            99,
            71,
            93,
            107,
            1,
            -68,
            -114,
            70,
            39,
            42,
            50,
            87,
            37,
            -41,
            56,
            0,
            15,
            106,
            123,
            -56,
            -86,
            8,
            64,
            -107,
            92,
            0,
            48,
            118,
            -46,
            -45,
            37,
            -114,
            19,
            99,
            58,
            -27,
            69,
            45,
            -2,
            -1,
            71,
            -99,
            78,
            -115,
            -86,
            -7,
            -72,
            78,
            -76,
            20,
            -85,
            -106,
            -115,
            -97,
            -126,
            -96,
            26,
            -46,
            122,
            -38,
            107,
            120,
            -70,
            111,
            127,
            -13,
            -43,
            86,
            -125,
            -92,
            22,
            -101,
            51,
            4,
            48,
            -17,
            109,
            -13,
            -61,
            -66,
            41,
            2,
            0,
            0,
            -112,
            -115,
            -102,
            -101,
            58,
            -71,
            0,
            -64,
            9,
            -64,
            -41,
            116,
            -20,
            23,
            -23,
            -19,
            -14,
            34,
            -54,
            74,
            71,
            46,
            -119,
            -3,
            -109,
            -98,
            115,
            -53,
            -114,
            -34,
            -97,
            -21,
            108,
            -64,
            -86,
            35,
            108,
            -13,
            -120,
            44,
            61,
            -17,
            -25,
            -39,
            10,
            -97,
            -13,
            -7,
            65,
            122,
            -18,
            -17,
            -79,
            53,
            -1,
            39,
            79,
            11,
            -120,
            -12,
            18,
            15,
            13,
            48,
            92,
            126,
            116,
            -34,
            -28,
            22,
            73,
            54,
            -70,
            -123,
            -8,
            49,
            -50,
            56,
            -43,
            -84,
            115,
            -125,
            84,
            95,
            -74,
            86,
            10,
            12,
            48,
            30,
            80,
            -83,
            -67,
            -21,
            -5,
            -39,
            -52,
            7,
            0,
            80,
            -77,
            -80,
            -115,
            -29,
            -28,
            -10,
            -6,
            121,
            -94,
            92,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            -32,
            7,
            96,
            43,
            -27,
            99,
            29,
            -67,
            59,
            -50,
            -4,
            105,
            48,
            8,
            -86,
            -120,
            114,
            -21,
            -82,
            35,
            16,
            8,
            4,
            2,
            -127,
            -88,
            28,
            -65,
            108,
            -7,
            -73,
            85,
            66,
            -36,
            22,
            -27,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "daa97664-b256-4ce5-a82f-9faa353871ef",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "4189a92c-812b-4f84-b7fd-566eb4487e75",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Peking",
        "lastUpdate": 1448099237816,
        "uniqueIdentifier": "03bd7084-7b9c-48d8-b5ce-eab2a32f01c4",
        "description": "Peking Logistics Centre"
      },
      {
        "location": {
          "continent": "Asia",
          "country": {
            "isoNumber3": 392,
            "name": "Japan",
            "isoAlpha2": "JP",
            "isoAlpha3": "JPN"
          },
          "state": null,
          "town": "Tokio",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            1,
            -106,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -103,
            49,
            78,
            -61,
            64,
            16,
            69,
            7,
            46,
            2,
            2,
            33,
            81,
            -92,
            -96,
            -128,
            36,
            -126,
            -96,
            -72,
            33,
            -95,
            9,
            78,
            -55,
            49,
            114,
            -125,
            -8,
            70,
            57,
            -126,
            83,
            32,
            74,
            -96,
            -95,
            68,
            -71,
            66,
            42,
            58,
            52,
            -20,
            40,
            88,
            32,
            107,
            109,
            111,
            -52,
            38,
            -69,
            107,
            -1,
            47,
            -3,
            46,
            -2,
            51,
            -13,
            36,
            -17,
            -114,
            21,
            34,
            8,
            -126,
            32,
            8,
            -126,
            -96,
            31,
            -11,
            -58,
            49,
            23,
            56,
            21,
            119,
            71,
            -15,
            -94,
            59,
            122,
            -104,
            -117,
            123,
            -29,
            73,
            124,
            117,
            55,
            25,
            110,
            60,
            -67,
            -40,
            87,
            -113,
            82,
            43,
            -85,
            43,
            61,
            100,
            -3,
            72,
            111,
            89,
            -97,
            69,
            115,
            84,
            -122,
            -85,
            -96,
            101,
            9,
            -124,
            109,
            -100,
            -2,
            -11,
            111,
            -109,
            102,
            -50,
            63,
            111,
            -93,
            39,
            -103,
            -51,
            -120,
            -80,
            69,
            8,
            -34,
            -40,
            120,
            120,
            -47,
            -27,
            -3,
            52,
            106,
            26,
            0,
            -103,
            -55,
            -42,
            89,
            16,
            -92,
            -1,
            125,
            -16,
            -16,
            45,
            113,
            72,
            -74,
            126,
            -14,
            -86,
            -48,
            117,
            64,
            0,
            -42,
            59,
            -71,
            126,
            120,
            64,
            111,
            -34,
            15,
            63,
            -96,
            -27,
            -50,
            -18,
            95,
            21,
            30,
            121,
            15,
            -32,
            -102,
            -10,
            -74,
            -113,
            -48,
            71,
            -121,
            -72,
            -60,
            73,
            -99,
            -61,
            -75,
            -96,
            78,
            82,
            86,
            -53,
            -39,
            -42,
            8,
            0,
            109,
            7,
            32,
            90,
            28,
            29,
            114,
            -34,
            79,
            39,
            52,
            51,
            -39,
            47,
            -8,
            125,
            99,
            -109,
            -5,
            90,
            50,
            117,
            -75,
            -100,
            127,
            60,
            -75,
            30,
            -64,
            -13,
            -39,
            1,
            -25,
            -3,
            114,
            74,
            -113,
            -74,
            1,
            72,
            -90,
            -82,
            -106,
            115,
            0,
            -70,
            119,
            114,
            -43,
            -95,
            -56,
            54,
            0,
            -55,
            -12,
            -18,
            -3,
            111,
            21,
            0,
            -18,
            -45,
            -79,
            90,
            52,
            -122,
            -66,
            3,
            -112,
            30,
            -91,
            87,
            103,
            91,
            -32,
            103,
            -97,
            -8,
            -21,
            -122,
            94,
            -43,
            -17,
            83,
            -27,
            121,
            -34,
            85,
            0,
            116,
            -49,
            72,
            -106,
            100,
            74,
            -74,
            -31,
            58,
            28,
            57,
            3,
            80,
            -27,
            74,
            0,
            118,
            -66,
            7,
            -62,
            0,
            -96,
            51,
            0,
            0,
            -128,
            -89,
            0,
            108,
            109,
            -126,
            117,
            -43,
            -104,
            85,
            -72,
            113,
            0,
            -74,
            -35,
            3,
            -22,
            -86,
            49,
            -101,
            32,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            4,
            15,
            32,
            -55,
            123,
            117,
            110,
            -1,
            -49,
            73,
            -55,
            -44,
            -43,
            34,
            8,
            -126,
            32,
            8,
            -126,
            32,
            -88,
            -98,
            -66,
            1,
            -78,
            -100,
            -118,
            63,
            -15,
            32,
            -87,
            -113,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "b3f51bf1-11ac-4037-bc20-8f03320e5a88",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "9c8f0641-3369-48dd-be84-7845d9c720ae",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Tokio",
        "lastUpdate": 1448099264285,
        "uniqueIdentifier": "ba8565ff-9186-4a9c-9b31-60ed9267133b",
        "description": "Tokio Logistics Centre"
      },
      {
        "location": {
          "continent": "Asia",
          "country": {
            "isoNumber3": 682,
            "name": "Saudi Arabia",
            "isoAlpha2": "SA",
            "isoAlpha3": "SAU"
          },
          "state": null,
          "town": "Abu Dhabi",
          "postcode": null,
          "street": null,
          "housenumber": null,
          "position": null
        },
        "icon": {
          "data": [
            -119,
            80,
            78,
            71,
            13,
            10,
            26,
            10,
            0,
            0,
            0,
            13,
            73,
            72,
            68,
            82,
            0,
            0,
            0,
            64,
            0,
            0,
            0,
            64,
            8,
            6,
            0,
            0,
            0,
            -86,
            105,
            113,
            -34,
            0,
            0,
            2,
            -114,
            73,
            68,
            65,
            84,
            120,
            -38,
            -19,
            -105,
            79,
            75,
            27,
            65,
            24,
            -58,
            -13,
            17,
            -4,
            8,
            -126,
            -121,
            -126,
            23,
            -67,
            121,
            106,
            -119,
            39,
            5,
            -5,
            5,
            60,
            88,
            68,
            61,
            40,
            109,
            122,
            -86,
            55,
            73,
            54,
            17,
            76,
            -76,
            21,
            -1,
            -128,
            1,
            69,
            27,
            91,
            115,
            80,
            15,
            -58,
            -118,
            -12,
            80,
            11,
            -46,
            -117,
            120,
            40,
            88,
            122,
            -23,
            81,
            63,
            -126,
            -33,
            96,
            -100,
            119,
            113,
            100,
            93,
            -9,
            -35,
            -35,
            -103,
            -99,
            -75,
            -101,
            -16,
            -68,
            -16,
            -64,
            50,
            -69,
            51,
            -17,
            -13,
            -2,
            -26,
            79,
            38,
            -71,
            28,
            2,
            -127,
            64,
            32,
            16,
            8,
            68,
            68,
            52,
            -86,
            78,
            126,
            -73,
            86,
            -70,
            -2,
            82,
            43,
            -119,
            -58,
            -118,
            -45,
            -107,
            57,
            127,
            -46,
            19,
            121,
            35,
            -113,
            -28,
            -43,
            122,
            2,
            26,
            92,
            -55,
            77,
            -78,
            -28,
            -12,
            39,
            54,
            45,
            -57,
            -112,
            102,
            -69,
            109,
            -116,
            -93,
            38,
            71,
            -55,
            98,
            -31,
            -59,
            85,
            -17,
            -64,
            94,
            -103,
            -102,
            -105,
            102,
            27,
            -2,
            -79,
            -88,
            -51,
            112,
            101,
            118,
            115,
            -2,
            -56,
            -69,
            -43,
            -103,
            15,
            72,
            112,
            -84,
            61,
            -34,
            98,
            -79,
            -60,
            -114,
            39,
            -33,
            25,
            76,
            -48,
            113,
            -104,
            -57,
            -108,
            1,
            -60,
            79,
            32,
            103,
            -72,
            21,
            53,
            -106,
            103,
            53,
            -76,
            -98,
            -37,
            31,
            -97,
            -96,
            90,
            -68,
            -31,
            6,
            -1,
            90,
            117,
            -58,
            19,
            -51,
            120,
            -108,
            98,
            -84,
            8,
            -14,
            -64,
            -10,
            -105,
            -34,
            115,
            54,
            14,
            24,
            83,
            -70,
            -22,
            100,
            78,
            -94,
            56,
            -65,
            56,
            108,
            95,
            11,
            7,
            117,
            -82,
            -16,
            122,
            80,
            -80,
            26,
            -55,
            95,
            -121,
            44,
            -7,
            -85,
            -92,
            -59,
            123,
            -74,
            -60,
            21,
            -105,
            -25,
            -35,
            -56,
            -32,
            109,
            -104,
            -57,
            116,
            1,
            48,
            9,
            -62,
            79,
            102,
            -69,
            43,
            -63,
            -60,
            -97,
            -55,
            57,
            -32,
            -60,
            -35,
            2,
            114,
            -74,
            -50,
            109,
            23,
            31,
            117,
            56,
            50,
            -5,
            -33,
            -79,
            119,
            23,
            -48,
            0,
            -112,
            86,
            -15,
            -38,
            57,
            -1,
            7,
            0,
            -7,
            -35,
            110,
            -38,
            0,
            -126,
            46,
            55,
            -39,
            1,
            -112,
            122,
            -15,
            26,
            121,
            1,
            0,
            0,
            0,
            0,
            0,
            0,
            -32,
            -103,
            1,
            -48,
            109,
            -19,
            104,
            107,
            93,
            68,
            -23,
            -37,
            78,
            -3,
            79,
            -112,
            -30,
            -12,
            13,
            -70,
            17,
            102,
            -22,
            34,
            -12,
            -17,
            -9,
            -91,
            72,
            83,
            -103,
            -65,
            9,
            2,
            -64,
            -67,
            -47,
            -51,
            -123,
            -110,
            24,
            -53,
            15,
            -72,
            -94,
            103,
            -43,
            -82,
            -38,
            72,
            97,
            109,
            92,
            127,
            0,
            0,
            0,
            -100,
            1,
            0,
            0,
            0,
            -19,
            14,
            -32,
            -17,
            -59,
            47,
            113,
            -78,
            -77,
            33,
            -106,
            -33,
            79,
            -70,
            -94,
            103,
            106,
            -53,
            20,
            -128,
            -77,
            -125,
            61,
            -25,
            -25,
            97,
            83,
            -24,
            42,
            -86,
            -128,
            -26,
            -57,
            -7,
            -121,
            -62,
            -3,
            -94,
            119,
            81,
            -3,
            77,
            60,
            81,
            45,
            -103,
            0,
            112,
            -7,
            -29,
            -108,
            45,
            94,
            -119,
            -66,
            -23,
            72,
            0,
            81,
            -123,
            -5,
            -43,
            81,
            0,
            -50,
            -113,
            -10,
            -75,
            1,
            80,
            -97,
            -114,
            0,
            -80,
            -65,
            -74,
            -88,
            93,
            -68,
            18,
            -11,
            109,
            123,
            0,
            -90,
            -59,
            115,
            91,
            33,
            19,
            0,
            -66,
            -17,
            109,
            -57,
            7,
            80,
            -104,
            96,
            85,
            -103,
            26,
            117,
            21,
            -10,
            77,
            92,
            0,
            97,
            -98,
            -84,
            2,
            40,
            79,
            -113,
            -117,
            -55,
            -95,
            -105,
            98,
            125,
            -18,
            67,
            -94,
            21,
            80,
            -101,
            121,
            35,
            94,
            -67,
            -24,
            113,
            69,
            -49,
            73,
            86,
            -64,
            -89,
            -39,
            -126,
            -21,
            -119,
            -68,
            -91,
            6,
            -128,
            -110,
            120,
            -1,
            -76,
            -112,
            40,
            -23,
            65,
            125,
            69,
            27,
            -128,
            42,
            -36,
            47,
            93,
            0,
            -108,
            -101,
            60,
            -8,
            125,
            -111,
            87,
            -85,
            0,
            90,
            -37,
            -11,
            39,
            73,
            -68,
            -46,
            1,
            48,
            -44,
            -41,
            -53,
            2,
            24,
            -18,
            -17,
            -43,
            2,
            16,
            -26,
            -119,
            60,
            91,
            3,
            -16,
            -71,
            86,
            -74,
            6,
            -128,
            43,
            -98,
            91,
            5,
            -90,
            0,
            -56,
            -77,
            53,
            0,
            -107,
            -73,
            19,
            109,
            7,
            -128,
            60,
            91,
            3,
            16,
            -76,
            -1,
            -77,
            14,
            -64,
            123,
            14,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            0,
            2,
            -127,
            64,
            32,
            16,
            8,
            -60,
            -93,
            -72,
            3,
            35,
            -101,
            105,
            32,
            70,
            30,
            -121,
            115,
            0,
            0,
            0,
            0,
            73,
            69,
            78,
            68,
            -82,
            66,
            96,
            -126
          ],
          "imageType": "png"
        },
        "next": null,
        "procedures": [
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Unload",
            "lastUpdate": 0,
            "uniqueIdentifier": "145a66e0-0087-4f71-a4d8-4c0330633726",
            "description": null
          },
          {
            "category": "Costs not accounted",
            "cost": {
              "Min": 500.0,
              "Max": 500.0
            },
            "time": {
              "Min": 60.0,
              "Max": 60.0
            },
            "timeType": "MINUTES",
            "cotwo": {
              "Min": 100.0,
              "Max": 100.0
            },
            "id": "#-1:-1",
            "name": "Load",
            "lastUpdate": 0,
            "uniqueIdentifier": "293cf57e-cde9-4d12-afd3-767a2de7d817",
            "description": null
          }
        ],
        "events": [],
        "id": null,
        "name": "Abu Dhabi",
        "lastUpdate": 1448099359735,
        "uniqueIdentifier": "0f413e8f-acc3-4bb0-b883-b94e85b5273b",
        "description": "Abu Dhabi Logistics Centre"
      }
    ],
    "basicProcedures": [
      {
        "category": "CheckUp",
        "cost": {
          "Min": 20.0,
          "Max": 20.0
        },
        "time": {
          "Min": 1.0,
          "Max": 1.0
        },
        "timeType": "HOURS",
        "cotwo": {
          "Min": 0.0,
          "Max": 0.0
        },
        "id": null,
        "name": "CheckUp",
        "lastUpdate": 1448100609375,
        "uniqueIdentifier": "e1128862-f0de-43ec-b554-5462ddbe4be3",
        "description": null
      },
      {
        "category": "Costs not accounted",
        "cost": {
          "Min": 500.0,
          "Max": 500.0
        },
        "time": {
          "Min": 3.0,
          "Max": 3.0
        },
        "timeType": "HOURS",
        "cotwo": {
          "Min": 50.0,
          "Max": 50.0
        },
        "id": null,
        "name": "Unload",
        "lastUpdate": 1448100642245,
        "uniqueIdentifier": "3690d36a-0a4a-44b0-8a6a-533e7e9d90bd",
        "description": null
      },
      {
        "category": "Load",
        "cost": {
          "Min": 500.0,
          "Max": 500.0
        },
        "time": {
          "Min": 3.0,
          "Max": 3.0
        },
        "timeType": "HOURS",
        "cotwo": {
          "Min": 50.0,
          "Max": 50.0
        },
        "id": null,
        "name": "Load",
        "lastUpdate": 1448100694362,
        "uniqueIdentifier": "f817ae0d-783c-4071-a70d-4ae0a76baa4d",
        "description": null
      }
    ]
  }
]